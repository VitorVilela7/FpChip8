library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity c8_prog_rom is
   port( CLK      : in std_logic;
         ADDR     : in natural range 0 to 21331;
         Q        : out std_logic_vector(7 downto 0));
end c8_prog_rom;

architecture rtl of c8_prog_rom is
   type rom_t is array (natural range <>) of std_logic_vector(7 downto 0);
   
   signal program : rom_t(0 to 21075) := (
		x"00", x"E0", x"6C", x"00", x"4C", x"00", x"6E", x"0F", x"A2", x"03", x"60", x"20", x"F0", x"55", x"00", x"E0",
		x"22", x"BE", x"22", x"76", x"22", x"8E", x"22", x"5E", x"22", x"46", x"12", x"10", x"61", x"00", x"62", x"17",
		x"63", x"04", x"41", x"10", x"00", x"EE", x"A2", x"E8", x"F1", x"1E", x"F0", x"65", x"40", x"00", x"12", x"34",
		x"F0", x"29", x"D2", x"35", x"71", x"01", x"72", x"05", x"64", x"03", x"84", x"12", x"34", x"00", x"12", x"22",
		x"62", x"17", x"73", x"06", x"12", x"22", x"64", x"03", x"84", x"E2", x"65", x"03", x"85", x"D2", x"94", x"50",
		x"00", x"EE", x"44", x"03", x"00", x"EE", x"64", x"01", x"84", x"E4", x"22", x"A6", x"12", x"46", x"64", x"03",
		x"84", x"E2", x"65", x"03", x"85", x"D2", x"94", x"50", x"00", x"EE", x"44", x"00", x"00", x"EE", x"64", x"FF",
		x"84", x"E4", x"22", x"A6", x"12", x"5E", x"64", x"0C", x"84", x"E2", x"65", x"0C", x"85", x"D2", x"94", x"50",
		x"00", x"EE", x"44", x"00", x"00", x"EE", x"64", x"FC", x"84", x"E4", x"22", x"A6", x"12", x"76", x"64", x"0C",
		x"84", x"E2", x"65", x"0C", x"85", x"D2", x"94", x"50", x"00", x"EE", x"44", x"0C", x"00", x"EE", x"64", x"04",
		x"84", x"E4", x"22", x"A6", x"12", x"8E", x"A2", x"E8", x"F4", x"1E", x"F0", x"65", x"A2", x"E8", x"FE", x"1E",
		x"F0", x"55", x"60", x"00", x"A2", x"E8", x"F4", x"1E", x"F0", x"55", x"8E", x"40", x"00", x"EE", x"3C", x"00",
		x"12", x"D2", x"22", x"1C", x"22", x"D8", x"22", x"1C", x"A2", x"F8", x"FD", x"1E", x"F0", x"65", x"8D", x"00",
		x"00", x"EE", x"7C", x"FF", x"CD", x"0F", x"00", x"EE", x"7D", x"01", x"60", x"0F", x"8D", x"02", x"ED", x"9E",
		x"12", x"D8", x"ED", x"A1", x"12", x"E2", x"00", x"EE", x"01", x"02", x"03", x"04", x"05", x"06", x"07", x"08",
		x"09", x"0A", x"0B", x"0C", x"0D", x"0E", x"0F", x"00", x"0D", x"00", x"01", x"02", x"04", x"05", x"06", x"08",
		x"09", x"0A", x"0C", x"0E", x"03", x"07", x"0B", x"0F", x"84", x"E4", x"22", x"A6", x"12", x"76", x"64", x"0C",
		x"84", x"E2", x"65", x"0C", x"85", x"D2", x"94", x"50", x"00", x"EE", x"44", x"0C", x"00", x"EE", x"64", x"04",
		x"84", x"E4", x"22", x"A6", x"12", x"8E", x"A2", x"E8", x"F4", x"1E", x"F0", x"65", x"A2", x"E8", x"FE", x"1E",
		x"F0", x"55", x"60", x"00", x"A2", x"E8", x"F4", x"1E", x"F0", x"55", x"8E", x"40", x"00", x"EE", x"3C", x"00",
		x"12", x"D2", x"22", x"1C", x"22", x"D8", x"22", x"1C", x"A2", x"F8", x"FD", x"1E", x"F0", x"65", x"8D", x"00",
		x"00", x"EE", x"7C", x"FF", x"CD", x"0F", x"00", x"EE", x"7D", x"01", x"60", x"0F", x"8D", x"02", x"ED", x"9E",
		x"12", x"D8", x"ED", x"A1", x"12", x"E2", x"00", x"EE", x"01", x"02", x"03", x"04", x"05", x"06", x"07", x"08",
		x"09", x"0A", x"0B", x"0C", x"0D", x"0E", x"0F", x"00", x"0D", x"00", x"01", x"02", x"04", x"05", x"06", x"08",
		x"12", x"1A", x"32", x"2E", x"30", x"30", x"20", x"43", x"2E", x"20", x"45", x"67", x"65", x"62", x"65", x"72",
		x"67", x"20", x"31", x"38", x"2F", x"38", x"2D", x"27", x"39", x"31", x"80", x"03", x"81", x"13", x"A8", x"C8",
		x"F1", x"55", x"60", x"05", x"A8", x"CC", x"F0", x"55", x"87", x"73", x"86", x"63", x"27", x"72", x"00", x"E0",
		x"27", x"94", x"6E", x"40", x"87", x"E2", x"6E", x"27", x"87", x"E1", x"68", x"1A", x"69", x"0C", x"6A", x"38",
		x"6B", x"00", x"6C", x"02", x"6D", x"1A", x"27", x"50", x"A8", x"ED", x"DA", x"B4", x"DC", x"D4", x"23", x"D0",
		x"3E", x"00", x"12", x"7C", x"A8", x"CC", x"F0", x"65", x"85", x"00", x"C4", x"FF", x"84", x"52", x"24", x"F6",
		x"C4", x"FF", x"84", x"52", x"26", x"1E", x"60", x"01", x"E0", x"A1", x"27", x"D6", x"36", x"F7", x"12", x"4E",
		x"8E", x"60", x"28", x"7A", x"6E", x"64", x"28", x"7A", x"27", x"D6", x"12", x"2A", x"F0", x"07", x"40", x"00",
		x"13", x"10", x"80", x"80", x"80", x"06", x"81", x"A0", x"81", x"06", x"80", x"15", x"40", x"00", x"12", x"9A",
		x"40", x"01", x"12", x"9A", x"40", x"FF", x"12", x"9A", x"12", x"C8", x"80", x"90", x"80", x"06", x"81", x"B0",
		x"81", x"06", x"80", x"15", x"40", x"00", x"12", x"B2", x"40", x"01", x"12", x"B2", x"40", x"FF", x"12", x"B2",
		x"12", x"C8", x"A8", x"ED", x"DA", x"B4", x"6A", x"38", x"6B", x"00", x"DA", x"B4", x"6E", x"F3", x"87", x"E2",
		x"6E", x"04", x"87", x"E1", x"6E", x"32", x"28", x"7A", x"80", x"80", x"80", x"06", x"81", x"C0", x"81", x"06",
		x"80", x"15", x"40", x"00", x"12", x"E0", x"40", x"01", x"12", x"E0", x"40", x"FF", x"12", x"E0", x"12", x"54",
		x"80", x"90", x"80", x"06", x"81", x"D0", x"81", x"06", x"80", x"15", x"40", x"00", x"12", x"F8", x"40", x"01",
		x"12", x"F8", x"40", x"FF", x"12", x"F8", x"12", x"54", x"A8", x"ED", x"DC", x"D4", x"6C", x"02", x"6D", x"1A",
		x"DC", x"D4", x"6E", x"CF", x"87", x"E2", x"6E", x"20", x"87", x"E1", x"6E", x"19", x"28", x"7A", x"12", x"54",
		x"60", x"3F", x"28", x"A8", x"27", x"50", x"A8", x"ED", x"DA", x"B4", x"DC", x"D4", x"6E", x"40", x"87", x"E3",
		x"80", x"70", x"80", x"E2", x"30", x"00", x"12", x"32", x"8E", x"60", x"28", x"7A", x"28", x"8A", x"00", x"E0",
		x"66", x"11", x"67", x"0A", x"A8", x"CA", x"27", x"E6", x"66", x"11", x"67", x"10", x"A8", x"C8", x"27", x"E6",
		x"64", x"00", x"65", x"08", x"66", x"00", x"67", x"0F", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69",
		x"60", x"03", x"28", x"A8", x"3E", x"00", x"13", x"C6", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69",
		x"74", x"02", x"75", x"02", x"34", x"30", x"13", x"48", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69",
		x"60", x"03", x"28", x"A8", x"3E", x"00", x"13", x"C6", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69",
		x"76", x"02", x"36", x"16", x"13", x"68", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69", x"60", x"03",
		x"28", x"A8", x"3E", x"00", x"13", x"C6", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69", x"74", x"FE",
		x"75", x"FE", x"34", x"00", x"13", x"86", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69", x"60", x"03",
		x"28", x"A8", x"3E", x"00", x"13", x"C6", x"AB", x"19", x"D4", x"69", x"AB", x"22", x"D5", x"69", x"76", x"FE",
		x"36", x"00", x"13", x"A6", x"13", x"48", x"AB", x"22", x"D5", x"69", x"AB", x"2B", x"D5", x"69", x"12", x"1A",
		x"83", x"70", x"6E", x"03", x"83", x"E2", x"84", x"80", x"85", x"90", x"6E", x"06", x"EE", x"A1", x"14", x"32",
		x"6E", x"03", x"EE", x"A1", x"14", x"4A", x"6E", x"08", x"EE", x"A1", x"14", x"62", x"6E", x"07", x"EE", x"A1",
		x"14", x"7A", x"43", x"03", x"75", x"02", x"43", x"00", x"75", x"FE", x"43", x"02", x"74", x"02", x"43", x"01",
		x"74", x"FE", x"80", x"40", x"81", x"50", x"27", x"BA", x"82", x"00", x"6E", x"08", x"80", x"E2", x"30", x"00",
		x"14", x"92", x"6E", x"07", x"80", x"20", x"82", x"E2", x"42", x"05", x"14", x"9A", x"42", x"06", x"14", x"B2",
		x"42", x"07", x"14", x"EC", x"27", x"50", x"6E", x"FC", x"87", x"E2", x"87", x"31", x"88", x"40", x"89", x"50",
		x"17", x"50", x"80", x"40", x"81", x"50", x"71", x"02", x"27", x"BA", x"82", x"00", x"6E", x"08", x"80", x"E2",
		x"30", x"00", x"13", x"F2", x"63", x"03", x"75", x"02", x"14", x"0E", x"80", x"40", x"81", x"50", x"71", x"FE",
		x"27", x"BA", x"82", x"00", x"6E", x"08", x"80", x"E2", x"30", x"00", x"13", x"F2", x"63", x"00", x"75", x"FE",
		x"14", x"0E", x"80", x"40", x"81", x"50", x"70", x"02", x"27", x"BA", x"82", x"00", x"6E", x"08", x"80", x"E2",
		x"30", x"00", x"13", x"F2", x"63", x"02", x"74", x"02", x"14", x"0E", x"80", x"40", x"81", x"50", x"70", x"FE",
		x"27", x"BA", x"82", x"00", x"6E", x"08", x"80", x"E2", x"30", x"00", x"13", x"F2", x"63", x"01", x"74", x"FE",
		x"14", x"0E", x"27", x"50", x"D8", x"94", x"8E", x"F0", x"00", x"EE", x"6E", x"F0", x"80", x"E2", x"80", x"31",
		x"F0", x"55", x"A8", x"F1", x"D4", x"54", x"76", x"01", x"61", x"05", x"F0", x"07", x"40", x"00", x"F1", x"18",
		x"14", x"24", x"6E", x"F0", x"80", x"E2", x"80", x"31", x"F0", x"55", x"A8", x"F5", x"D4", x"54", x"76", x"04",
		x"80", x"A0", x"81", x"B0", x"27", x"BA", x"6E", x"F0", x"80", x"E2", x"30", x"00", x"14", x"D2", x"6E", x"0C",
		x"87", x"E3", x"80", x"C0", x"81", x"D0", x"27", x"BA", x"6E", x"F0", x"80", x"E2", x"30", x"00", x"14", x"E4",
		x"6E", x"30", x"87", x"E3", x"60", x"FF", x"F0", x"18", x"F0", x"15", x"14", x"24", x"43", x"01", x"64", x"3A",
		x"43", x"02", x"64", x"00", x"14", x"24", x"82", x"70", x"83", x"70", x"6E", x"0C", x"82", x"E2", x"80", x"A0",
		x"81", x"B0", x"27", x"BA", x"A8", x"ED", x"6E", x"F0", x"80", x"E2", x"30", x"00", x"15", x"24", x"DA", x"B4",
		x"42", x"0C", x"7B", x"02", x"42", x"00", x"7B", x"FE", x"42", x"08", x"7A", x"02", x"42", x"04", x"7A", x"FE",
		x"DA", x"B4", x"00", x"EE", x"6E", x"80", x"F1", x"07", x"31", x"00", x"15", x"D4", x"34", x"00", x"15", x"D4",
		x"81", x"00", x"83", x"0E", x"3F", x"00", x"15", x"56", x"83", x"90", x"83", x"B5", x"4F", x"00", x"15", x"8C",
		x"33", x"00", x"15", x"74", x"87", x"E3", x"83", x"80", x"83", x"A5", x"4F", x"00", x"15", x"BC", x"33", x"00",
		x"15", x"A4", x"87", x"E3", x"15", x"D4", x"83", x"80", x"83", x"A5", x"4F", x"00", x"15", x"BC", x"33", x"00",
		x"15", x"A4", x"87", x"E3", x"83", x"90", x"83", x"B5", x"4F", x"00", x"15", x"8C", x"33", x"00", x"15", x"74",
		x"87", x"E3", x"15", x"D4", x"63", x"40", x"81", x"32", x"41", x"00", x"15", x"D4", x"DA", x"B4", x"7B", x"02",
		x"DA", x"B4", x"6E", x"F3", x"87", x"E2", x"62", x"0C", x"87", x"21", x"00", x"EE", x"63", x"10", x"81", x"32",
		x"41", x"00", x"15", x"D4", x"DA", x"B4", x"7B", x"FE", x"DA", x"B4", x"6E", x"F3", x"87", x"E2", x"62", x"00",
		x"87", x"21", x"00", x"EE", x"63", x"20", x"81", x"32", x"41", x"00", x"15", x"D4", x"DA", x"B4", x"7A", x"02",
		x"DA", x"B4", x"6E", x"F3", x"87", x"E2", x"62", x"08", x"87", x"21", x"00", x"EE", x"63", x"80", x"81", x"32",
		x"41", x"00", x"15", x"D4", x"DA", x"B4", x"7A", x"FE", x"DA", x"B4", x"6E", x"F3", x"87", x"E2", x"62", x"04",
		x"87", x"21", x"00", x"EE", x"C1", x"F0", x"80", x"12", x"30", x"00", x"15", x"E4", x"6E", x"0C", x"87", x"E3",
		x"82", x"E3", x"15", x"0E", x"DA", x"B4", x"80", x"0E", x"4F", x"00", x"15", x"F2", x"62", x"04", x"7A", x"FE",
		x"16", x"14", x"80", x"0E", x"4F", x"00", x"15", x"FE", x"62", x"0C", x"7B", x"02", x"16", x"14", x"80", x"0E",
		x"4F", x"00", x"16", x"0A", x"62", x"08", x"7A", x"02", x"16", x"14", x"80", x"0E", x"4F", x"00", x"15", x"DC",
		x"62", x"00", x"7B", x"FE", x"DA", x"B4", x"6E", x"F3", x"87", x"E2", x"87", x"21", x"00", x"EE", x"82", x"70",
		x"83", x"70", x"6E", x"30", x"82", x"E2", x"80", x"C0", x"81", x"D0", x"27", x"BA", x"A8", x"ED", x"6E", x"F0",
		x"80", x"E2", x"30", x"00", x"16", x"4C", x"DC", x"D4", x"42", x"30", x"7D", x"02", x"42", x"00", x"7D", x"FE",
		x"42", x"20", x"7C", x"02", x"42", x"10", x"7C", x"FE", x"DC", x"D4", x"00", x"EE", x"6E", x"80", x"F1", x"07",
		x"31", x"00", x"17", x"04", x"34", x"00", x"17", x"04", x"81", x"00", x"83", x"0E", x"4F", x"00", x"16", x"7E",
		x"83", x"90", x"83", x"D5", x"4F", x"00", x"16", x"B6", x"33", x"00", x"16", x"9C", x"87", x"E3", x"83", x"80",
		x"83", x"C5", x"4F", x"00", x"16", x"EA", x"33", x"00", x"16", x"D0", x"87", x"E3", x"17", x"04", x"83", x"80",
		x"83", x"C5", x"4F", x"00", x"16", x"EA", x"33", x"00", x"16", x"D0", x"87", x"E3", x"83", x"90", x"83", x"D5",
		x"4F", x"00", x"16", x"B6", x"33", x"00", x"16", x"9C", x"87", x"E3", x"17", x"04", x"63", x"40", x"81", x"32",
		x"41", x"00", x"17", x"04", x"DC", x"D4", x"7D", x"02", x"DC", x"D4", x"87", x"E3", x"6E", x"CF", x"87", x"E2",
		x"62", x"30", x"87", x"21", x"00", x"EE", x"63", x"10", x"81", x"32", x"41", x"00", x"17", x"04", x"DC", x"D4",
		x"7D", x"FE", x"DC", x"D4", x"87", x"E3", x"6E", x"CF", x"87", x"E2", x"62", x"00", x"87", x"21", x"00", x"EE",
		x"63", x"20", x"81", x"32", x"41", x"00", x"17", x"04", x"DC", x"D4", x"7C", x"02", x"DC", x"D4", x"87", x"E3",
		x"6E", x"CF", x"87", x"E2", x"62", x"20", x"87", x"21", x"00", x"EE", x"63", x"80", x"81", x"32", x"41", x"00",
		x"17", x"04", x"DC", x"D4", x"7C", x"FE", x"DC", x"D4", x"87", x"E3", x"6E", x"CF", x"87", x"E2", x"62", x"10",
		x"87", x"21", x"00", x"EE", x"C1", x"F0", x"80", x"12", x"30", x"00", x"17", x"16", x"87", x"E3", x"6E", x"30",
		x"87", x"E3", x"82", x"E3", x"16", x"36", x"DC", x"D4", x"80", x"0E", x"4F", x"00", x"17", x"24", x"62", x"90",
		x"7C", x"FE", x"17", x"46", x"80", x"0E", x"4F", x"00", x"17", x"30", x"62", x"30", x"7D", x"02", x"17", x"46",
		x"80", x"0E", x"4F", x"00", x"17", x"3C", x"62", x"A0", x"7C", x"02", x"17", x"46", x"80", x"0E", x"4F", x"00",
		x"17", x"0C", x"62", x"00", x"7D", x"FE", x"DC", x"D4", x"6E", x"4F", x"87", x"E2", x"87", x"21", x"00", x"EE",
		x"80", x"70", x"6E", x"03", x"80", x"E2", x"80", x"0E", x"81", x"80", x"81", x"94", x"6E", x"02", x"81", x"E2",
		x"41", x"00", x"70", x"01", x"80", x"0E", x"80", x"0E", x"A8", x"CD", x"F0", x"1E", x"D8", x"94", x"8E", x"F0",
		x"00", x"EE", x"6E", x"00", x"A9", x"19", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"F3", x"65",
		x"AB", x"34", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"F3", x"55", x"7E", x"01", x"3E", x"80",
		x"17", x"74", x"00", x"EE", x"82", x"23", x"83", x"33", x"6E", x"0F", x"80", x"20", x"81", x"30", x"27", x"BE",
		x"80", x"E2", x"80", x"0E", x"A8", x"F9", x"F0", x"1E", x"D2", x"32", x"72", x"02", x"32", x"40", x"17", x"9A",
		x"82", x"23", x"73", x"02", x"43", x"20", x"00", x"EE", x"17", x"9A", x"70", x"02", x"71", x"02", x"80", x"06",
		x"81", x"06", x"81", x"0E", x"81", x"0E", x"81", x"0E", x"81", x"0E", x"AB", x"34", x"F1", x"1E", x"F1", x"1E",
		x"F0", x"1E", x"F0", x"65", x"00", x"EE", x"A8", x"CC", x"F0", x"65", x"80", x"06", x"F0", x"55", x"60", x"01",
		x"E0", x"A1", x"17", x"E0", x"00", x"EE", x"F1", x"65", x"6E", x"01", x"84", x"43", x"82", x"00", x"83", x"10",
		x"65", x"10", x"83", x"55", x"4F", x"00", x"82", x"E5", x"4F", x"00", x"18", x"0C", x"65", x"27", x"82", x"55",
		x"4F", x"00", x"18", x"0C", x"80", x"20", x"81", x"30", x"84", x"E4", x"17", x"F0", x"F4", x"29", x"D6", x"75",
		x"76", x"06", x"84", x"43", x"82", x"00", x"83", x"10", x"65", x"E8", x"83", x"55", x"4F", x"00", x"82", x"E5",
		x"4F", x"00", x"18", x"34", x"65", x"03", x"82", x"55", x"4F", x"00", x"18", x"34", x"80", x"20", x"81", x"30",
		x"84", x"E4", x"18", x"18", x"F4", x"29", x"D6", x"75", x"76", x"06", x"84", x"43", x"82", x"00", x"83", x"10",
		x"65", x"64", x"83", x"55", x"4F", x"00", x"82", x"E5", x"4F", x"00", x"18", x"54", x"80", x"20", x"81", x"30",
		x"84", x"E4", x"18", x"40", x"F4", x"29", x"D6", x"75", x"76", x"06", x"84", x"43", x"82", x"00", x"83", x"10",
		x"65", x"0A", x"83", x"55", x"4F", x"00", x"18", x"6E", x"81", x"30", x"84", x"E4", x"18", x"60", x"F4", x"29",
		x"D6", x"75", x"76", x"06", x"F1", x"29", x"D6", x"75", x"00", x"EE", x"A8", x"C8", x"F1", x"65", x"81", x"E4",
		x"3F", x"00", x"70", x"01", x"A8", x"C8", x"F1", x"55", x"00", x"EE", x"A8", x"C8", x"F3", x"65", x"8E", x"00",
		x"8E", x"25", x"4F", x"00", x"00", x"EE", x"3E", x"00", x"18", x"A2", x"8E", x"10", x"8E", x"35", x"4F", x"00",
		x"00", x"EE", x"A8", x"CA", x"F1", x"55", x"00", x"EE", x"8E", x"E3", x"62", x"0F", x"63", x"FF", x"61", x"10",
		x"E2", x"A1", x"18", x"C4", x"81", x"34", x"31", x"00", x"18", x"B0", x"61", x"10", x"80", x"34", x"30", x"00",
		x"18", x"B0", x"00", x"EE", x"6E", x"01", x"00", x"EE", x"00", x"00", x"00", x"00", x"05", x"00", x"50", x"70",
		x"20", x"00", x"50", x"70", x"20", x"00", x"60", x"30", x"60", x"00", x"60", x"30", x"60", x"00", x"30", x"60",
		x"30", x"00", x"30", x"60", x"30", x"00", x"20", x"70", x"50", x"00", x"20", x"70", x"50", x"00", x"20", x"70",
		x"70", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"80", x"00", x"00", x"00", x"00", x"00", x"C0", x"00", x"00", x"00", x"80", x"80", x"00",
		x"00", x"C0", x"80", x"80", x"80", x"C0", x"00", x"80", x"00", x"0C", x"08", x"08", x"08", x"08", x"08", x"08",
		x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0D", x"0C", x"08", x"08", x"08", x"08", x"08", x"08",
		x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0D", x"0A", x"65", x"05", x"05", x"05", x"05", x"E5",
		x"05", x"05", x"E5", x"05", x"05", x"05", x"05", x"C5", x"0A", x"0A", x"65", x"05", x"05", x"05", x"05", x"E5",
		x"05", x"05", x"E5", x"05", x"05", x"05", x"05", x"C5", x"0A", x"0A", x"05", x"0C", x"08", x"08", x"0F", x"05",
		x"0C", x"0D", x"05", x"08", x"08", x"08", x"0D", x"05", x"0E", x"0F", x"05", x"0C", x"08", x"08", x"0F", x"05",
		x"0C", x"0D", x"05", x"08", x"08", x"08", x"0D", x"05", x"0A", x"0A", x"05", x"0A", x"65", x"06", x"05", x"95",
		x"0A", x"0A", x"35", x"05", x"05", x"C5", x"0A", x"35", x"05", x"05", x"95", x"0A", x"65", x"05", x"05", x"95",
		x"0A", x"0A", x"35", x"05", x"06", x"C5", x"0A", x"05", x"0A", x"0A", x"05", x"0F", x"05", x"08", x"08", x"08",
		x"08", x"08", x"0C", x"08", x"0F", x"05", x"08", x"08", x"08", x"08", x"08", x"0F", x"05", x"08", x"08", x"0C",
		x"08", x"08", x"08", x"08", x"0F", x"05", x"0F", x"05", x"0A", x"0A", x"75", x"05", x"B5", x"05", x"05", x"05",
		x"05", x"C5", x"0A", x"65", x"05", x"B5", x"05", x"E5", x"05", x"05", x"E5", x"05", x"B5", x"05", x"C5", x"0A",
		x"65", x"05", x"05", x"05", x"05", x"B5", x"05", x"D5", x"0A", x"0A", x"05", x"0C", x"08", x"08", x"08", x"08",
		x"0D", x"05", x"0F", x"05", x"0C", x"08", x"0F", x"05", x"08", x"0F", x"05", x"08", x"08", x"0D", x"05", x"0F",
		x"05", x"0C", x"08", x"08", x"08", x"08", x"0D", x"05", x"0A", x"0F", x"05", x"0F", x"65", x"05", x"05", x"C5",
		x"0A", x"35", x"E5", x"95", x"0A", x"65", x"05", x"B0", x"05", x"05", x"B5", x"05", x"C5", x"0A", x"35", x"E5",
		x"95", x"0A", x"65", x"05", x"05", x"C5", x"0F", x"05", x"0F", x"07", x"74", x"05", x"D5", x"08", x"0F", x"05",
		x"0E", x"0F", x"05", x"08", x"0F", x"05", x"0C", x"08", x"08", x"08", x"08", x"0D", x"05", x"08", x"0F", x"05",
		x"08", x"0F", x"05", x"08", x"0F", x"75", x"05", x"D4", x"07", x"0A", x"05", x"0A", x"35", x"05", x"05", x"F5",
		x"05", x"05", x"B5", x"05", x"05", x"D5", x"08", x"08", x"0D", x"0C", x"08", x"0F", x"75", x"05", x"05", x"B5",
		x"05", x"05", x"F5", x"05", x"05", x"95", x"0A", x"05", x"0A", x"0A", x"05", x"08", x"08", x"08", x"0D", x"05",
		x"0C", x"08", x"08", x"08", x"0D", x"35", x"05", x"C5", x"0A", x"0A", x"65", x"05", x"95", x"0C", x"08", x"08",
		x"08", x"0D", x"05", x"0C", x"08", x"08", x"0F", x"05", x"0A", x"0A", x"75", x"05", x"06", x"C5", x"0A", x"05",
		x"08", x"08", x"08", x"08", x"08", x"08", x"0F", x"05", x"08", x"0F", x"05", x"08", x"08", x"08", x"08", x"08",
		x"08", x"0F", x"05", x"0A", x"65", x"06", x"05", x"D5", x"0A", x"0A", x"05", x"0C", x"0D", x"05", x"0A", x"35",
		x"05", x"05", x"05", x"05", x"E5", x"05", x"05", x"F5", x"05", x"05", x"F5", x"05", x"05", x"E5", x"05", x"05",
		x"05", x"05", x"95", x"0A", x"05", x"0C", x"0D", x"05", x"0A", x"0A", x"05", x"08", x"0F", x"05", x"08", x"08",
		x"08", x"08", x"08", x"0F", x"05", x"0C", x"0D", x"05", x"08", x"0F", x"05", x"0C", x"0D", x"05", x"08", x"08",
		x"08", x"08", x"08", x"0F", x"05", x"08", x"0F", x"05", x"0A", x"0A", x"35", x"05", x"05", x"B5", x"05", x"05",
		x"05", x"05", x"05", x"05", x"95", x"0A", x"0A", x"35", x"05", x"05", x"95", x"0A", x"0A", x"35", x"05", x"05",
		x"05", x"05", x"05", x"05", x"B5", x"05", x"05", x"95", x"0A", x"08", x"08", x"08", x"08", x"08", x"08", x"08",
		x"08", x"08", x"08", x"08", x"08", x"0F", x"08", x"08", x"08", x"08", x"08", x"0F", x"08", x"08", x"08", x"08",
		x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0F", x"3C", x"42", x"99", x"99", x"42", x"3C", x"01",
		x"10", x"0F", x"78", x"84", x"32", x"32", x"84", x"78", x"00", x"10", x"E0", x"78", x"FC", x"FE", x"FE", x"84",
		x"78", x"00", x"10", x"E0", x"12", x"17", x"42", x"4C", x"49", x"54", x"5A", x"20", x"42", x"79", x"20", x"44",
		x"61", x"76", x"69", x"64", x"20", x"57", x"49", x"4E", x"54", x"45", x"52", x"A3", x"41", x"60", x"04", x"61",
		x"09", x"62", x"0E", x"67", x"04", x"D0", x"1E", x"F2", x"1E", x"70", x"0C", x"30", x"40", x"12", x"21", x"F0",
		x"0A", x"00", x"E0", x"22", x"D9", x"F0", x"0A", x"00", x"E0", x"8E", x"70", x"A3", x"1E", x"6B", x"1F", x"CC",
		x"1F", x"8C", x"C4", x"DC", x"B2", x"3F", x"01", x"12", x"49", x"DC", x"B2", x"12", x"39", x"CA", x"07", x"7A",
		x"01", x"7B", x"FE", x"DC", x"B2", x"7A", x"FF", x"3A", x"00", x"12", x"4D", x"7E", x"FF", x"3E", x"00", x"12",
		x"39", x"6B", x"00", x"8C", x"70", x"6D", x"00", x"6E", x"00", x"A3", x"1B", x"DD", x"E3", x"3F", x"00", x"12",
		x"C1", x"3B", x"00", x"12", x"81", x"60", x"05", x"E0", x"9E", x"12", x"87", x"6B", x"01", x"88", x"D0", x"78",
		x"02", x"89", x"E0", x"79", x"03", x"A3", x"1E", x"D8", x"91", x"81", x"F0", x"60", x"05", x"F0", x"15", x"F0",
		x"07", x"30", x"00", x"12", x"8B", x"3B", x"01", x"12", x"AB", x"A3", x"1E", x"31", x"01", x"D8", x"91", x"79",
		x"01", x"39", x"20", x"12", x"AB", x"6B", x"00", x"31", x"00", x"7C", x"FF", x"4C", x"00", x"12", x"BB", x"A3",
		x"1B", x"DD", x"E3", x"7D", x"02", x"3D", x"40", x"12", x"B9", x"6D", x"00", x"7E", x"01", x"12", x"65", x"00",
		x"E0", x"77", x"02", x"12", x"2D", x"A3", x"1B", x"DD", x"E3", x"60", x"14", x"61", x"02", x"62", x"0B", x"A3",
		x"20", x"D0", x"1B", x"F2", x"1E", x"70", x"08", x"30", x"2C", x"12", x"CD", x"12", x"D7", x"60", x"0A", x"61",
		x"0D", x"62", x"05", x"A3", x"07", x"D0", x"15", x"F2", x"1E", x"70", x"08", x"30", x"2A", x"12", x"E1", x"80",
		x"70", x"70", x"FE", x"80", x"06", x"A3", x"87", x"F0", x"33", x"F2", x"65", x"60", x"2D", x"F1", x"29", x"61",
		x"0D", x"D0", x"15", x"70", x"05", x"F2", x"29", x"D0", x"15", x"00", x"EE", x"83", x"82", x"83", x"82", x"FB",
		x"E8", x"08", x"88", x"05", x"E2", x"BE", x"A0", x"B8", x"20", x"3E", x"80", x"80", x"80", x"80", x"F8", x"80",
		x"F8", x"FC", x"C0", x"C0", x"F9", x"81", x"DB", x"CB", x"FB", x"00", x"FA", x"8A", x"9A", x"99", x"F8", x"EF",
		x"2A", x"E8", x"29", x"29", x"00", x"6F", x"68", x"2E", x"4C", x"8F", x"BE", x"A0", x"B8", x"B0", x"BE", x"00",
		x"BE", x"22", x"3E", x"34", x"B2", x"D8", x"D8", x"00", x"C3", x"C3", x"00", x"D8", x"D8", x"00", x"C3", x"C3",
		x"00", x"D8", x"D8", x"C0", x"C0", x"00", x"C0", x"C0", x"00", x"C0", x"C0", x"00", x"C0", x"C0", x"00", x"DB",
		x"DB", x"DB", x"DB", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"DB", x"DB", x"DB",
		x"DB", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"18", x"18", x"00", x"18", x"18", x"DB", x"DB", x"00",
		x"03", x"03", x"00", x"18", x"18", x"00", x"C0", x"C0", x"00", x"DB", x"DB", x"A2", x"5B", x"60", x"0B", x"61",
		x"03", x"62", x"07", x"D0", x"17", x"70", x"07", x"F2", x"1E", x"D0", x"17", x"70", x"07", x"F2", x"1E", x"D0",
		x"17", x"70", x"07", x"F2", x"1E", x"D0", x"17", x"70", x"07", x"F2", x"1E", x"D0", x"17", x"70", x"05", x"F2",
		x"1E", x"D0", x"17", x"F2", x"1E", x"A2", x"5A", x"C0", x"3F", x"C1", x"1F", x"62", x"01", x"63", x"01", x"D0",
		x"11", x"64", x"02", x"F4", x"15", x"F4", x"07", x"34", x"00", x"12", x"3A", x"D0", x"11", x"80", x"24", x"81",
		x"34", x"D0", x"11", x"41", x"00", x"63", x"01", x"41", x"1F", x"63", x"FF", x"40", x"00", x"62", x"01", x"40",
		x"3F", x"62", x"FF", x"12", x"36", x"80", x"78", x"CC", x"C0", x"C0", x"C0", x"CC", x"78", x"CC", x"CC", x"CC",
		x"FC", x"CC", x"CC", x"CC", x"FC", x"30", x"30", x"30", x"30", x"30", x"FC", x"F8", x"CC", x"CC", x"F8", x"C0",
		x"C0", x"C0", x"00", x"00", x"00", x"F0", x"00", x"00", x"00", x"78", x"CC", x"CC", x"78", x"CC", x"CC", x"78",
		x"6E", x"05", x"65", x"00", x"6B", x"06", x"6A", x"00", x"A3", x"0C", x"DA", x"B1", x"7A", x"04", x"3A", x"40",
		x"12", x"08", x"7B", x"02", x"3B", x"12", x"12", x"06", x"6C", x"20", x"6D", x"1F", x"A3", x"10", x"DC", x"D1",
		x"22", x"F6", x"60", x"00", x"61", x"00", x"A3", x"12", x"D0", x"11", x"70", x"08", x"A3", x"0E", x"D0", x"11",
		x"60", x"40", x"F0", x"15", x"F0", x"07", x"30", x"00", x"12", x"34", x"C6", x"0F", x"67", x"1E", x"68", x"01",
		x"69", x"FF", x"A3", x"0E", x"D6", x"71", x"A3", x"10", x"DC", x"D1", x"60", x"04", x"E0", x"A1", x"7C", x"FE",
		x"60", x"06", x"E0", x"A1", x"7C", x"02", x"60", x"3F", x"8C", x"02", x"DC", x"D1", x"A3", x"0E", x"D6", x"71",
		x"86", x"84", x"87", x"94", x"60", x"3F", x"86", x"02", x"61", x"1F", x"87", x"12", x"47", x"1F", x"12", x"AC",
		x"46", x"00", x"68", x"01", x"46", x"3F", x"68", x"FF", x"47", x"00", x"69", x"01", x"D6", x"71", x"3F", x"01",
		x"12", x"AA", x"47", x"1F", x"12", x"AA", x"60", x"05", x"80", x"75", x"3F", x"00", x"12", x"AA", x"60", x"01",
		x"F0", x"18", x"80", x"60", x"61", x"FC", x"80", x"12", x"A3", x"0C", x"D0", x"71", x"60", x"FE", x"89", x"03",
		x"22", x"F6", x"75", x"01", x"22", x"F6", x"45", x"60", x"12", x"DE", x"12", x"46", x"69", x"FF", x"80", x"60",
		x"80", x"C5", x"3F", x"01", x"12", x"CA", x"61", x"02", x"80", x"15", x"3F", x"01", x"12", x"E0", x"80", x"15",
		x"3F", x"01", x"12", x"EE", x"80", x"15", x"3F", x"01", x"12", x"E8", x"60", x"20", x"F0", x"18", x"A3", x"0E",
		x"7E", x"FF", x"80", x"E0", x"80", x"04", x"61", x"00", x"D0", x"11", x"3E", x"00", x"12", x"30", x"12", x"DE",
		x"78", x"FF", x"48", x"FE", x"68", x"FF", x"12", x"EE", x"78", x"01", x"48", x"02", x"68", x"01", x"60", x"04",
		x"F0", x"18", x"69", x"FF", x"12", x"70", x"A3", x"14", x"F5", x"33", x"F2", x"65", x"F1", x"29", x"63", x"37",
		x"64", x"00", x"D3", x"45", x"73", x"05", x"F2", x"29", x"D3", x"45", x"00", x"EE", x"E0", x"00", x"80", x"00",
		x"FC", x"00", x"AA", x"00", x"00", x"00", x"00", x"00", x"00", x"E0", x"64", x"00", x"65", x"00", x"A2", x"0A",
		x"12", x"0C", x"CC", x"33", x"66", x"1E", x"D4", x"52", x"D4", x"62", x"74", x"08", x"44", x"40", x"12", x"1A",
		x"12", x"0E", x"A2", x"1E", x"12", x"2C", x"FF", x"FF", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0", x"C0",
		x"C0", x"C0", x"FF", x"FF", x"64", x"0D", x"65", x"09", x"D4", x"5E", x"74", x"0A", x"A2", x"3A", x"D4", x"5E",
		x"12", x"48", x"FF", x"FF", x"C3", x"C3", x"C3", x"C3", x"C3", x"FF", x"FF", x"C3", x"C3", x"C3", x"C3", x"C3",
		x"74", x"0A", x"A2", x"50", x"D4", x"5E", x"12", x"5E", x"C3", x"C3", x"C3", x"C3", x"C3", x"66", x"66", x"66",
		x"66", x"66", x"3C", x"3C", x"18", x"18", x"74", x"0A", x"A2", x"66", x"D4", x"5E", x"12", x"74", x"FF", x"FF",
		x"C0", x"C0", x"C0", x"C0", x"FF", x"FF", x"C0", x"C0", x"C0", x"C0", x"FF", x"FF", x"6A", x"01", x"6B", x"04",
		x"6C", x"0E", x"6D", x"00", x"A2", x"81", x"12", x"A6", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
		x"FF", x"FF", x"00", x"E0", x"64", x"00", x"65", x"00", x"D4", x"58", x"74", x"08", x"44", x"40", x"22", x"9E",
		x"45", x"20", x"12", x"A4", x"12", x"90", x"64", x"00", x"75", x"08", x"00", x"EE", x"12", x"AE", x"60", x"0F",
		x"E0", x"9E", x"12", x"A8", x"12", x"8A", x"4A", x"01", x"22", x"D0", x"4A", x"02", x"23", x"8A", x"4A", x"03",
		x"23", x"B8", x"4A", x"04", x"23", x"E0", x"4A", x"05", x"24", x"18", x"4A", x"06", x"24", x"78", x"4A", x"07",
		x"24", x"E6", x"4A", x"08", x"25", x"10", x"13", x"18", x"A2", x"81", x"64", x"02", x"65", x"02", x"D4", x"58",
		x"65", x"0A", x"D4", x"58", x"65", x"12", x"D4", x"58", x"64", x"0A", x"65", x"05", x"D4", x"53", x"64", x"12",
		x"D4", x"53", x"64", x"1A", x"D4", x"53", x"64", x"22", x"D4", x"53", x"64", x"2A", x"D4", x"53", x"64", x"32",
		x"D4", x"53", x"A2", x"FE", x"13", x"0A", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC",
		x"FC", x"FC", x"75", x"03", x"74", x"02", x"D4", x"5C", x"74", x"06", x"75", x"09", x"D4", x"53", x"00", x"EE",
		x"A2", x"80", x"DB", x"C1", x"4F", x"01", x"13", x"72", x"60", x"02", x"E0", x"A1", x"6D", x"02", x"60", x"04",
		x"E0", x"A1", x"6D", x"04", x"60", x"06", x"E0", x"A1", x"6D", x"06", x"60", x"08", x"E0", x"A1", x"6D", x"08",
		x"DB", x"C1", x"4D", x"02", x"7C", x"FF", x"4D", x"04", x"7B", x"FF", x"4D", x"06", x"7B", x"01", x"4D", x"08",
		x"7C", x"01", x"4B", x"40", x"13", x"5E", x"4B", x"FF", x"13", x"64", x"60", x"02", x"F0", x"15", x"F0", x"07",
		x"30", x"00", x"13", x"56", x"13", x"18", x"7A", x"01", x"4A", x"09", x"15", x"3A", x"6B", x"01", x"A2", x"81",
		x"12", x"8A", x"7A", x"FF", x"6B", x"3E", x"A2", x"81", x"12", x"8A", x"60", x"03", x"F0", x"18", x"60", x"0F",
		x"E0", x"9E", x"13", x"78", x"6A", x"01", x"6B", x"04", x"6C", x"0E", x"6D", x"00", x"A2", x"81", x"00", x"E0",
		x"12", x"8A", x"64", x"00", x"65", x"11", x"A2", x"81", x"D4", x"53", x"74", x"08", x"D4", x"53", x"74", x"08",
		x"75", x"FF", x"D4", x"53", x"74", x"08", x"75", x"FF", x"D4", x"53", x"74", x"08", x"D4", x"53", x"74", x"08",
		x"D4", x"53", x"74", x"08", x"75", x"01", x"D4", x"53", x"74", x"08", x"75", x"01", x"D4", x"53", x"00", x"EE",
		x"64", x"00", x"65", x"11", x"A2", x"81", x"D4", x"53", x"74", x"08", x"D4", x"53", x"74", x"08", x"75", x"02",
		x"D4", x"52", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08",
		x"D4", x"51", x"74", x"08", x"D4", x"51", x"00", x"EE", x"64", x"00", x"65", x"13", x"A2", x"81", x"D4", x"51",
		x"A2", x"80", x"74", x"08", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"A2", x"81", x"D4", x"51",
		x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"52", x"74", x"08", x"75", x"FF", x"D4", x"53", x"74", x"08",
		x"D4", x"54", x"74", x"08", x"75", x"FF", x"D4", x"56", x"74", x"08", x"75", x"FF", x"D4", x"58", x"00", x"EE",
		x"64", x"00", x"65", x"12", x"A2", x"81", x"D4", x"58", x"74", x"08", x"D4", x"58", x"74", x"08", x"D4", x"58",
		x"74", x"08", x"D4", x"58", x"74", x"08", x"D4", x"58", x"74", x"08", x"D4", x"58", x"74", x"08", x"D4", x"58",
		x"A2", x"80", x"75", x"FF", x"74", x"20", x"D4", x"51", x"75", x"FF", x"D4", x"51", x"75", x"FF", x"D4", x"51",
		x"75", x"FF", x"D4", x"51", x"75", x"FF", x"D4", x"51", x"75", x"FF", x"D4", x"51", x"75", x"FF", x"D4", x"51",
		x"75", x"FF", x"D4", x"51", x"75", x"FF", x"A2", x"81", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08",
		x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"00", x"EE",
		x"64", x"00", x"65", x"09", x"A2", x"81", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51",
		x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"A2", x"80", x"75", x"01",
		x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01",
		x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01",
		x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01",
		x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01", x"D4", x"51", x"75", x"01",
		x"A2", x"81", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"00", x"EE", x"64", x"00",
		x"65", x"1A", x"A2", x"81", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08",
		x"D4", x"51", x"74", x"08", x"D4", x"51", x"75", x"FF", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08",
		x"D4", x"51", x"74", x"08", x"D4", x"51", x"00", x"EE", x"64", x"00", x"65", x"19", x"A2", x"81", x"D4", x"51",
		x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51",
		x"75", x"FF", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51", x"74", x"08", x"D4", x"51",
		x"00", x"EE", x"00", x"E0", x"67", x"03", x"68", x"03", x"A5", x"44", x"15", x"5C", x"AE", x"AA", x"EA", x"4A",
		x"4E", x"00", x"A4", x"A4", x"A4", x"A5", x"E2", x"00", x"5D", x"55", x"55", x"55", x"9D", x"00", x"C8", x"48",
		x"48", x"40", x"48", x"00", x"D7", x"85", x"A5", x"4A", x"77", x"08", x"D7", x"85", x"77", x"08", x"A5", x"50",
		x"D7", x"85", x"77", x"08", x"A5", x"56", x"D7", x"85", x"15", x"70", x"12", x"1A", x"43", x"4F", x"4E", x"4E",
		x"45", x"43", x"54", x"34", x"20", x"62", x"79", x"20", x"44", x"61", x"76", x"69", x"64", x"20", x"57", x"49",
		x"4E", x"54", x"45", x"52", x"A2", x"BB", x"F6", x"65", x"A2", x"B4", x"F6", x"55", x"69", x"00", x"68", x"01",
		x"6B", x"00", x"6D", x"0F", x"6E", x"1F", x"A2", x"A5", x"60", x"0D", x"61", x"32", x"62", x"00", x"D0", x"2F",
		x"D1", x"2F", x"72", x"0F", x"32", x"1E", x"12", x"34", x"D0", x"21", x"D1", x"21", x"72", x"01", x"60", x"0A",
		x"A2", x"9F", x"D0", x"21", x"D1", x"21", x"A2", x"9F", x"DD", x"E1", x"FC", x"0A", x"DD", x"E1", x"4C", x"05",
		x"12", x"7E", x"3C", x"04", x"12", x"6A", x"7B", x"FF", x"7D", x"FB", x"3D", x"0A", x"12", x"7A", x"6B", x"06",
		x"6D", x"2D", x"12", x"7A", x"3C", x"06", x"12", x"98", x"7B", x"01", x"7D", x"05", x"3D", x"32", x"12", x"7A",
		x"6B", x"00", x"6D", x"0F", x"DD", x"E1", x"12", x"50", x"A2", x"B4", x"FB", x"1E", x"F0", x"65", x"40", x"FC",
		x"12", x"98", x"8A", x"00", x"70", x"FB", x"F0", x"55", x"89", x"83", x"A2", x"9E", x"39", x"00", x"A2", x"A1",
		x"DD", x"A4", x"A2", x"9F", x"DD", x"E1", x"12", x"50", x"60", x"F0", x"F0", x"60", x"90", x"90", x"60", x"80",
		x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"1A", x"1A",
		x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"1A", x"6E", x"01", x"00", x"E0",
		x"6D", x"01", x"6A", x"01", x"6B", x"01", x"8C", x"D0", x"8C", x"E2", x"4C", x"00", x"12", x"20", x"88", x"D0",
		x"22", x"3E", x"3A", x"40", x"12", x"20", x"6A", x"01", x"7B", x"06", x"3C", x"3F", x"7D", x"01", x"3D", x"3F",
		x"12", x"0A", x"F0", x"0A", x"40", x"05", x"89", x"E4", x"8E", x"E4", x"3E", x"40", x"12", x"02", x"6A", x"1C",
		x"6B", x"0D", x"88", x"90", x"00", x"E0", x"22", x"3E", x"12", x"3C", x"A2", x"94", x"F8", x"33", x"F2", x"65",
		x"22", x"54", x"DA", x"B5", x"7A", x"04", x"81", x"20", x"22", x"54", x"DA", x"B5", x"7A", x"05", x"00", x"EE",
		x"83", x"10", x"83", x"34", x"83", x"34", x"83", x"14", x"A2", x"62", x"F3", x"1E", x"00", x"EE", x"E0", x"A0",
		x"A0", x"A0", x"E0", x"40", x"40", x"40", x"40", x"40", x"E0", x"20", x"E0", x"80", x"E0", x"E0", x"20", x"E0",
		x"20", x"E0", x"A0", x"A0", x"E0", x"20", x"20", x"E0", x"80", x"E0", x"20", x"E0", x"E0", x"80", x"E0", x"A0",
		x"E0", x"E0", x"20", x"20", x"20", x"20", x"E0", x"A0", x"E0", x"A0", x"E0", x"E0", x"A0", x"E0", x"20", x"E0",
		x"12", x"1D", x"48", x"49", x"44", x"44", x"45", x"4E", x"21", x"20", x"31", x"2E", x"30", x"20", x"42", x"79",
		x"20", x"44", x"61", x"76", x"69", x"64", x"20", x"57", x"49", x"4E", x"54", x"45", x"52", x"A4", x"3F", x"60",
		x"00", x"61", x"40", x"F1", x"55", x"A4", x"3F", x"60", x"00", x"F0", x"55", x"00", x"E0", x"A4", x"7E", x"60",
		x"0C", x"61", x"08", x"62", x"0F", x"D0", x"1F", x"70", x"08", x"F2", x"1E", x"30", x"34", x"12", x"35", x"F0",
		x"0A", x"00", x"E0", x"A4", x"C9", x"60", x"13", x"61", x"0D", x"62", x"04", x"D0", x"14", x"70", x"08", x"F2",
		x"1E", x"30", x"2B", x"12", x"4B", x"A4", x"1F", x"FF", x"65", x"A4", x"2F", x"FF", x"55", x"63", x"40", x"66",
		x"08", x"C1", x"0F", x"C2", x"0F", x"A4", x"2F", x"F1", x"1E", x"F0", x"65", x"84", x"00", x"A4", x"2F", x"F2",
		x"1E", x"F0", x"65", x"85", x"00", x"80", x"40", x"F0", x"55", x"A4", x"2F", x"F1", x"1E", x"80", x"50", x"F0",
		x"55", x"73", x"FF", x"33", x"00", x"12", x"61", x"00", x"E0", x"60", x"00", x"61", x"00", x"A4", x"77", x"D0",
		x"17", x"70", x"08", x"30", x"20", x"12", x"8F", x"60", x"00", x"71", x"08", x"31", x"20", x"12", x"8F", x"6C",
		x"00", x"6D", x"00", x"6E", x"00", x"A4", x"3F", x"F0", x"65", x"70", x"01", x"F0", x"55", x"23", x"B9", x"6A",
		x"10", x"23", x"5D", x"23", x"CD", x"8A", x"90", x"87", x"D0", x"88", x"E0", x"23", x"5D", x"23", x"CD", x"23",
		x"B9", x"A4", x"2F", x"F9", x"1E", x"F0", x"65", x"81", x"00", x"A4", x"2F", x"FA", x"1E", x"F0", x"65", x"50",
		x"10", x"13", x"2B", x"23", x"DF", x"60", x"20", x"24", x"01", x"23", x"DF", x"60", x"00", x"A4", x"2F", x"F9",
		x"1E", x"F0", x"55", x"A4", x"2F", x"FA", x"1E", x"F0", x"55", x"76", x"FF", x"36", x"00", x"12", x"A5", x"A4",
		x"3F", x"F1", x"65", x"82", x"00", x"80", x"15", x"3F", x"00", x"13", x"01", x"80", x"20", x"81", x"20", x"F1",
		x"55", x"00", x"E0", x"A5", x"19", x"60", x"10", x"61", x"07", x"62", x"0E", x"D0", x"1F", x"70", x"08", x"F2",
		x"1E", x"30", x"30", x"13", x"0B", x"A4", x"3F", x"F1", x"65", x"84", x"10", x"83", x"00", x"66", x"09", x"24",
		x"0B", x"66", x"0F", x"83", x"40", x"24", x"0B", x"F0", x"0A", x"12", x"25", x"23", x"DB", x"60", x"80", x"24",
		x"01", x"23", x"DB", x"A4", x"2F", x"FA", x"1E", x"F0", x"65", x"70", x"FF", x"23", x"F3", x"A4", x"41", x"F0",
		x"1E", x"D7", x"87", x"A4", x"77", x"D7", x"87", x"A4", x"2F", x"F9", x"1E", x"F0", x"65", x"70", x"FF", x"23",
		x"F3", x"A4", x"41", x"F0", x"1E", x"DD", x"E7", x"A4", x"77", x"DD", x"E7", x"12", x"A5", x"A4", x"71", x"DD",
		x"E7", x"FB", x"0A", x"DD", x"E7", x"3B", x"04", x"13", x"71", x"4D", x"00", x"13", x"5D", x"7D", x"F8", x"7C",
		x"FF", x"3B", x"06", x"13", x"7D", x"4D", x"18", x"13", x"5D", x"7D", x"08", x"7C", x"01", x"3B", x"02", x"13",
		x"89", x"4E", x"00", x"13", x"5D", x"7E", x"F8", x"7C", x"FC", x"3B", x"08", x"13", x"95", x"4E", x"18", x"13",
		x"5D", x"7E", x"08", x"7C", x"04", x"3B", x"05", x"13", x"5D", x"A4", x"2F", x"FC", x"1E", x"F0", x"65", x"40",
		x"00", x"13", x"5D", x"89", x"C0", x"99", x"A0", x"13", x"5D", x"70", x"FF", x"A4", x"77", x"DD", x"E7", x"A4",
		x"41", x"23", x"F3", x"F0", x"1E", x"DD", x"E7", x"00", x"EE", x"A4", x"D5", x"60", x"24", x"61", x"0A", x"62",
		x"0B", x"D0", x"1B", x"70", x"08", x"F2", x"1E", x"30", x"3C", x"13", x"C1", x"00", x"EE", x"60", x"34", x"61",
		x"10", x"A4", x"F1", x"D0", x"15", x"A4", x"F6", x"D0", x"15", x"00", x"EE", x"A4", x"FB", x"13", x"E1", x"A5",
		x"0A", x"60", x"24", x"61", x"0D", x"62", x"05", x"D0", x"15", x"70", x"08", x"F2", x"1E", x"30", x"3C", x"13",
		x"E7", x"00", x"EE", x"81", x"00", x"81", x"14", x"80", x"04", x"80", x"04", x"80", x"04", x"80", x"15", x"00",
		x"EE", x"F0", x"15", x"F0", x"07", x"30", x"00", x"14", x"03", x"00", x"EE", x"A4", x"2F", x"F3", x"33", x"F2",
		x"65", x"65", x"23", x"F1", x"29", x"D5", x"65", x"65", x"28", x"F2", x"29", x"D5", x"65", x"00", x"EE", x"01",
		x"02", x"03", x"04", x"08", x"07", x"06", x"05", x"05", x"06", x"07", x"08", x"04", x"03", x"02", x"01", x"01",
		x"02", x"03", x"04", x"08", x"07", x"06", x"05", x"05", x"06", x"07", x"08", x"04", x"03", x"02", x"01", x"00",
		x"00", x"FE", x"EE", x"C6", x"82", x"C6", x"EE", x"FE", x"FE", x"C6", x"C6", x"C6", x"FE", x"FE", x"C6", x"AA",
		x"82", x"AA", x"C6", x"FE", x"C6", x"82", x"82", x"82", x"C6", x"FE", x"BA", x"D6", x"EE", x"D6", x"BA", x"FE",
		x"EE", x"EE", x"82", x"EE", x"EE", x"FE", x"82", x"FE", x"82", x"FE", x"82", x"FE", x"AA", x"AA", x"AA", x"AA",
		x"AA", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"AA", x"D6", x"AA", x"D6", x"AA", x"FE", x"8B", x"88",
		x"F8", x"88", x"8B", x"00", x"00", x"00", x"00", x"00", x"F0", x"48", x"48", x"48", x"F2", x"EF", x"84", x"84",
		x"84", x"EF", x"00", x"08", x"08", x"0A", x"00", x"8A", x"8A", x"AA", x"AA", x"52", x"3C", x"92", x"92", x"92",
		x"3C", x"00", x"E2", x"A3", x"E3", x"00", x"8B", x"C8", x"A8", x"98", x"88", x"FA", x"83", x"E2", x"82", x"FA",
		x"00", x"28", x"B8", x"90", x"00", x"EF", x"88", x"8E", x"88", x"8F", x"21", x"21", x"A1", x"60", x"21", x"00",
		x"00", x"00", x"00", x"00", x"BC", x"22", x"3C", x"28", x"A4", x"89", x"8A", x"AB", x"52", x"97", x"51", x"D1",
		x"51", x"C0", x"00", x"00", x"15", x"6A", x"8A", x"8E", x"8A", x"6A", x"00", x"64", x"8A", x"8E", x"8A", x"6A",
		x"44", x"AA", x"AA", x"AA", x"44", x"00", x"CC", x"AA", x"CA", x"AA", x"AC", x"6E", x"88", x"4C", x"28", x"CE",
		x"00", x"04", x"0C", x"04", x"04", x"0E", x"0C", x"12", x"04", x"08", x"1E", x"63", x"94", x"94", x"94", x"63",
		x"38", x"A5", x"B8", x"A0", x"21", x"E1", x"01", x"C1", x"20", x"C1", x"89", x"8A", x"52", x"22", x"21", x"CF",
		x"28", x"2F", x"28", x"C8", x"02", x"82", x"02", x"00", x"02", x"FF", x"80", x"8F", x"90", x"8E", x"81", x"9E",
		x"80", x"91", x"91", x"9F", x"91", x"91", x"80", x"FF", x"00", x"3C", x"40", x"40", x"40", x"3C", x"00", x"7C",
		x"10", x"10", x"10", x"7C", x"00", x"FF", x"00", x"00", x"80", x"00", x"80", x"00", x"00", x"00", x"80", x"00",
		x"80", x"00", x"00", x"FF", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"01",
		x"01", x"FF", x"00", x"E0", x"A2", x"2A", x"60", x"0C", x"61", x"08", x"D0", x"1F", x"70", x"09", x"A2", x"39",
		x"D0", x"1F", x"A2", x"48", x"70", x"08", x"D0", x"1F", x"70", x"04", x"A2", x"57", x"D0", x"1F", x"70", x"08",
		x"A2", x"66", x"D0", x"1F", x"70", x"08", x"A2", x"75", x"D0", x"1F", x"12", x"28", x"FF", x"00", x"FF", x"00",
		x"3C", x"00", x"3C", x"00", x"3C", x"00", x"3C", x"00", x"FF", x"00", x"FF", x"FF", x"00", x"FF", x"00", x"38",
		x"00", x"3F", x"00", x"3F", x"00", x"38", x"00", x"FF", x"00", x"FF", x"80", x"00", x"E0", x"00", x"E0", x"00",
		x"80", x"00", x"80", x"00", x"E0", x"00", x"E0", x"00", x"80", x"F8", x"00", x"FC", x"00", x"3E", x"00", x"3F",
		x"00", x"3B", x"00", x"39", x"00", x"F8", x"00", x"F8", x"03", x"00", x"07", x"00", x"0F", x"00", x"BF", x"00",
		x"FB", x"00", x"F3", x"00", x"E3", x"00", x"43", x"E0", x"00", x"E0", x"00", x"80", x"00", x"80", x"00", x"80",
		x"00", x"80", x"00", x"E0", x"00", x"E0", x"12", x"25", x"53", x"50", x"41", x"43", x"45", x"20", x"49", x"4E",
		x"56", x"41", x"44", x"45", x"52", x"53", x"20", x"76", x"30", x"2E", x"39", x"20", x"42", x"79", x"20", x"44",
		x"61", x"76", x"69", x"64", x"20", x"57", x"49", x"4E", x"54", x"45", x"52", x"60", x"00", x"61", x"00", x"62",
		x"08", x"A3", x"D3", x"D0", x"18", x"71", x"08", x"F2", x"1E", x"31", x"20", x"12", x"2D", x"70", x"08", x"61",
		x"00", x"30", x"40", x"12", x"2D", x"69", x"05", x"6C", x"15", x"6E", x"00", x"23", x"87", x"60", x"0A", x"F0",
		x"15", x"F0", x"07", x"30", x"00", x"12", x"4B", x"23", x"87", x"7E", x"01", x"12", x"45", x"66", x"00", x"68",
		x"1C", x"69", x"00", x"6A", x"04", x"6B", x"0A", x"6C", x"04", x"6D", x"3C", x"6E", x"0F", x"00", x"E0", x"23",
		x"6B", x"23", x"47", x"FD", x"15", x"60", x"04", x"E0", x"9E", x"12", x"7D", x"23", x"6B", x"38", x"00", x"78",
		x"FF", x"23", x"6B", x"60", x"06", x"E0", x"9E", x"12", x"8B", x"23", x"6B", x"38", x"39", x"78", x"01", x"23",
		x"6B", x"36", x"00", x"12", x"9F", x"60", x"05", x"E0", x"9E", x"12", x"E9", x"66", x"01", x"65", x"1B", x"84",
		x"80", x"A3", x"CF", x"D4", x"51", x"A3", x"CF", x"D4", x"51", x"75", x"FF", x"35", x"FF", x"12", x"AD", x"66",
		x"00", x"12", x"E9", x"D4", x"51", x"3F", x"01", x"12", x"E9", x"D4", x"51", x"66", x"00", x"83", x"40", x"73",
		x"03", x"83", x"B5", x"62", x"F8", x"83", x"22", x"62", x"08", x"33", x"00", x"12", x"C9", x"23", x"73", x"82",
		x"06", x"43", x"08", x"12", x"D3", x"33", x"10", x"12", x"D5", x"23", x"73", x"82", x"06", x"33", x"18", x"12",
		x"DD", x"23", x"73", x"82", x"06", x"43", x"20", x"12", x"E7", x"33", x"28", x"12", x"E9", x"23", x"73", x"3E",
		x"00", x"13", x"07", x"79", x"06", x"49", x"18", x"69", x"00", x"6A", x"04", x"6B", x"0A", x"6C", x"04", x"7D",
		x"F4", x"6E", x"0F", x"00", x"E0", x"23", x"47", x"23", x"6B", x"FD", x"15", x"12", x"6F", x"F7", x"07", x"37",
		x"00", x"12", x"6F", x"FD", x"15", x"23", x"47", x"8B", x"A4", x"3B", x"12", x"13", x"1B", x"7C", x"02", x"6A",
		x"FC", x"3B", x"02", x"13", x"23", x"7C", x"02", x"6A", x"04", x"23", x"47", x"3C", x"18", x"12", x"6F", x"00",
		x"E0", x"A4", x"D3", x"60", x"14", x"61", x"08", x"62", x"0F", x"D0", x"1F", x"70", x"08", x"F2", x"1E", x"30",
		x"2C", x"13", x"33", x"F0", x"0A", x"00", x"E0", x"A6", x"F4", x"FE", x"65", x"12", x"25", x"A3", x"B7", x"F9",
		x"1E", x"61", x"08", x"23", x"5F", x"81", x"06", x"23", x"5F", x"81", x"06", x"23", x"5F", x"81", x"06", x"23",
		x"5F", x"7B", x"D0", x"00", x"EE", x"80", x"E0", x"80", x"12", x"30", x"00", x"DB", x"C6", x"7B", x"0C", x"00",
		x"EE", x"A3", x"CF", x"60", x"1C", x"D8", x"04", x"00", x"EE", x"23", x"47", x"8E", x"23", x"23", x"47", x"60",
		x"05", x"F0", x"18", x"F0", x"15", x"F0", x"07", x"30", x"00", x"13", x"7F", x"00", x"EE", x"6A", x"00", x"8D",
		x"E0", x"6B", x"04", x"E9", x"A1", x"12", x"57", x"A6", x"02", x"FD", x"1E", x"F0", x"65", x"30", x"FF", x"13",
		x"A5", x"6A", x"00", x"6B", x"04", x"6D", x"01", x"6E", x"01", x"13", x"8D", x"A5", x"00", x"F0", x"1E", x"DB",
		x"C6", x"7B", x"08", x"7D", x"01", x"7A", x"01", x"3A", x"07", x"13", x"8D", x"00", x"EE", x"3C", x"7E", x"FF",
		x"FF", x"99", x"99", x"7E", x"FF", x"FF", x"24", x"24", x"E7", x"7E", x"FF", x"3C", x"3C", x"7E", x"DB", x"81",
		x"42", x"3C", x"7E", x"FF", x"DB", x"10", x"38", x"7C", x"FE", x"00", x"00", x"7F", x"00", x"3F", x"00", x"7F",
		x"00", x"00", x"00", x"01", x"01", x"01", x"03", x"03", x"03", x"03", x"00", x"00", x"3F", x"20", x"20", x"20",
		x"20", x"20", x"20", x"20", x"20", x"3F", x"08", x"08", x"FF", x"00", x"00", x"FE", x"00", x"FC", x"00", x"FE",
		x"00", x"00", x"00", x"7E", x"42", x"42", x"62", x"62", x"62", x"62", x"00", x"00", x"FF", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"7D", x"00", x"41", x"7D", x"05", x"7D",
		x"7D", x"00", x"00", x"C2", x"C2", x"C6", x"44", x"6C", x"28", x"38", x"00", x"00", x"FF", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"F7", x"10", x"14", x"F7", x"F7", x"04",
		x"04", x"00", x"00", x"7C", x"44", x"FE", x"C2", x"C2", x"C2", x"C2", x"00", x"00", x"FF", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"EF", x"20", x"28", x"E8", x"E8", x"2F",
		x"2F", x"00", x"00", x"F9", x"85", x"C5", x"C5", x"C5", x"C5", x"F9", x"00", x"00", x"FF", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"BE", x"00", x"20", x"30", x"20", x"BE",
		x"BE", x"00", x"00", x"F7", x"04", x"E7", x"85", x"85", x"84", x"F4", x"00", x"00", x"FF", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"7F", x"00", x"3F", x"00", x"7F",
		x"00", x"00", x"00", x"EF", x"28", x"EF", x"00", x"E0", x"60", x"6F", x"00", x"00", x"FF", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"FF", x"00", x"00", x"FE", x"00", x"FC", x"00", x"FE",
		x"00", x"00", x"00", x"C0", x"00", x"C0", x"C0", x"C0", x"C0", x"C0", x"00", x"00", x"FC", x"04", x"04", x"04",
		x"04", x"04", x"04", x"04", x"04", x"FC", x"10", x"10", x"FF", x"F9", x"81", x"B9", x"8B", x"9A", x"9A", x"FA",
		x"00", x"FA", x"8A", x"9A", x"9A", x"9B", x"99", x"F8", x"E6", x"25", x"25", x"F4", x"34", x"34", x"34", x"00",
		x"17", x"14", x"34", x"37", x"36", x"26", x"C7", x"DF", x"50", x"50", x"5C", x"D8", x"D8", x"DF", x"00", x"DF",
		x"11", x"1F", x"12", x"1B", x"19", x"D9", x"7C", x"44", x"FE", x"86", x"86", x"86", x"FC", x"84", x"FE", x"82",
		x"82", x"FE", x"FE", x"80", x"C0", x"C0", x"C0", x"FE", x"FC", x"82", x"C2", x"C2", x"C2", x"FC", x"FE", x"80",
		x"F8", x"C0", x"C0", x"FE", x"FE", x"80", x"F0", x"C0", x"C0", x"C0", x"FE", x"80", x"BE", x"86", x"86", x"FE",
		x"86", x"86", x"FE", x"86", x"86", x"86", x"10", x"10", x"10", x"10", x"10", x"10", x"18", x"18", x"18", x"48",
		x"48", x"78", x"9C", x"90", x"B0", x"C0", x"B0", x"9C", x"80", x"80", x"C0", x"C0", x"C0", x"FE", x"EE", x"92",
		x"92", x"86", x"86", x"86", x"FE", x"82", x"86", x"86", x"86", x"86", x"7C", x"82", x"86", x"86", x"86", x"7C",
		x"FE", x"82", x"FE", x"C0", x"C0", x"C0", x"7C", x"82", x"C2", x"CA", x"C4", x"7A", x"FE", x"86", x"FE", x"90",
		x"9C", x"84", x"FE", x"C0", x"FE", x"02", x"02", x"FE", x"FE", x"10", x"30", x"30", x"30", x"30", x"82", x"82",
		x"C2", x"C2", x"C2", x"FE", x"82", x"82", x"82", x"EE", x"38", x"10", x"86", x"86", x"96", x"92", x"92", x"EE",
		x"82", x"44", x"38", x"38", x"44", x"82", x"82", x"82", x"FE", x"30", x"30", x"30", x"FE", x"02", x"1E", x"F0",
		x"80", x"FE", x"00", x"00", x"00", x"00", x"06", x"06", x"00", x"00", x"00", x"60", x"60", x"C0", x"00", x"00",
		x"00", x"00", x"00", x"00", x"18", x"18", x"18", x"18", x"00", x"18", x"7C", x"C6", x"0C", x"18", x"00", x"18",
		x"00", x"00", x"FE", x"FE", x"00", x"00", x"FE", x"82", x"86", x"86", x"86", x"FE", x"08", x"08", x"08", x"18",
		x"18", x"18", x"FE", x"02", x"FE", x"C0", x"C0", x"FE", x"FE", x"02", x"1E", x"06", x"06", x"FE", x"84", x"C4",
		x"C4", x"FE", x"04", x"04", x"FE", x"80", x"FE", x"06", x"06", x"FE", x"C0", x"C0", x"C0", x"FE", x"82", x"FE",
		x"FE", x"02", x"02", x"06", x"06", x"06", x"7C", x"44", x"FE", x"86", x"86", x"FE", x"FE", x"82", x"FE", x"06",
		x"06", x"06", x"44", x"FE", x"44", x"44", x"FE", x"44", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"6C",
		x"5A", x"00", x"0C", x"18", x"A8", x"30", x"4E", x"7E", x"00", x"12", x"18", x"66", x"6C", x"A8", x"5A", x"66",
		x"54", x"24", x"66", x"00", x"48", x"48", x"18", x"12", x"A8", x"06", x"90", x"A8", x"12", x"00", x"7E", x"30",
		x"12", x"A8", x"84", x"30", x"4E", x"72", x"18", x"66", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"90", x"54",
		x"78", x"A8", x"48", x"78", x"6C", x"72", x"A8", x"12", x"18", x"6C", x"72", x"66", x"54", x"90", x"A8", x"72",
		x"2A", x"18", x"A8", x"30", x"4E", x"7E", x"00", x"12", x"18", x"66", x"6C", x"A8", x"72", x"54", x"A8", x"5A",
		x"66", x"18", x"7E", x"18", x"4E", x"72", x"A8", x"72", x"2A", x"18", x"30", x"66", x"A8", x"30", x"4E", x"7E",
		x"00", x"6C", x"30", x"54", x"4E", x"9C", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"48", x"54", x"7E",
		x"18", x"A8", x"90", x"54", x"78", x"66", x"A8", x"6C", x"2A", x"30", x"5A", x"A8", x"84", x"30", x"72", x"2A",
		x"A8", x"D8", x"A8", x"00", x"4E", x"12", x"A8", x"E4", x"A2", x"A8", x"00", x"4E", x"12", x"A8", x"6C", x"2A",
		x"54", x"54", x"72", x"A8", x"84", x"30", x"72", x"2A", x"A8", x"DE", x"9C", x"A8", x"72", x"2A", x"18", x"A8",
		x"0C", x"54", x"48", x"5A", x"78", x"72", x"18", x"66", x"A8", x"72", x"18", x"42", x"42", x"6C", x"A8", x"72",
		x"2A", x"00", x"72", x"A8", x"72", x"2A", x"18", x"A8", x"30", x"4E", x"7E", x"00", x"12", x"18", x"66", x"6C",
		x"A8", x"30", x"4E", x"0C", x"66", x"18", x"00", x"6C", x"18", x"A8", x"72", x"2A", x"18", x"30", x"66", x"A8",
		x"1E", x"54", x"66", x"0C", x"18", x"9C", x"A8", x"24", x"54", x"54", x"12", x"A8", x"42", x"78", x"0C", x"3C",
		x"A8", x"AE", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"FF", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"00", x"63", x"80", x"61", x"1F", x"62",
		x"0F", x"22", x"32", x"A2", x"00", x"F3", x"1E", x"F0", x"0A", x"F0", x"55", x"40", x"00", x"12", x"1C", x"73",
		x"01", x"33", x"00", x"12", x"08", x"63", x"80", x"A2", x"00", x"F3", x"1E", x"F0", x"65", x"40", x"00", x"12",
		x"1C", x"73", x"01", x"43", x"00", x"12", x"1C", x"22", x"32", x"12", x"1E", x"40", x"02", x"72", x"FF", x"40",
		x"04", x"71", x"FF", x"40", x"06", x"71", x"01", x"40", x"08", x"72", x"01", x"A2", x"77", x"6A", x"E0", x"8A",
		x"12", x"6B", x"1F", x"81", x"B2", x"3A", x"00", x"72", x"01", x"6A", x"F0", x"8A", x"22", x"6B", x"0F", x"82",
		x"B2", x"3A", x"00", x"71", x"01", x"6B", x"1F", x"81", x"B2", x"D1", x"21", x"8A", x"10", x"6B", x"1F", x"8B",
		x"25", x"DA", x"B1", x"6A", x"3F", x"8A", x"15", x"DA", x"B1", x"8B", x"20", x"DA", x"B1", x"00", x"EE", x"01",
		x"80", x"12", x"4E", x"08", x"19", x"01", x"01", x"08", x"01", x"0F", x"01", x"01", x"09", x"08", x"09", x"0F",
		x"09", x"01", x"11", x"08", x"11", x"0F", x"11", x"01", x"19", x"0F", x"19", x"16", x"01", x"16", x"09", x"16",
		x"11", x"16", x"19", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"FC", x"00", x"A2", x"02", x"82", x"0E", x"F2",
		x"1E", x"82", x"06", x"F1", x"65", x"00", x"EE", x"A2", x"02", x"82", x"0E", x"F2", x"1E", x"82", x"06", x"F1",
		x"55", x"00", x"EE", x"6F", x"10", x"FF", x"15", x"FF", x"07", x"3F", x"00", x"12", x"46", x"00", x"EE", x"00",
		x"E0", x"62", x"00", x"22", x"2A", x"F2", x"29", x"D0", x"15", x"70", x"FF", x"71", x"FF", x"22", x"36", x"72",
		x"01", x"32", x"10", x"12", x"52", x"F2", x"0A", x"22", x"2A", x"A2", x"22", x"D0", x"17", x"22", x"42", x"D0",
		x"17", x"12", x"64", x"60", x"00", x"61", x"00", x"A2", x"22", x"C2", x"01", x"32", x"01", x"A2", x"1E", x"D0",
		x"14", x"70", x"04", x"30", x"40", x"12", x"04", x"60", x"00", x"71", x"04", x"31", x"20", x"12", x"04", x"12",
		x"1C", x"80", x"40", x"20", x"10", x"20", x"40", x"80", x"10", x"12", x"19", x"20", x"4D", x"45", x"52", x"4C",
		x"49", x"4E", x"20", x"42", x"79", x"20", x"44", x"61", x"76", x"69", x"64", x"20", x"57", x"49", x"4E", x"54",
		x"45", x"52", x"22", x"F9", x"A3", x"1D", x"60", x"10", x"61", x"00", x"22", x"CB", x"A3", x"31", x"60", x"0B",
		x"61", x"1B", x"22", x"CB", x"64", x"04", x"22", x"DF", x"65", x"00", x"62", x"28", x"22", x"C1", x"C2", x"03",
		x"80", x"20", x"A3", x"59", x"F5", x"1E", x"F0", x"55", x"60", x"17", x"61", x"08", x"63", x"01", x"83", x"22",
		x"33", x"00", x"70", x"0A", x"63", x"02", x"83", x"22", x"33", x"00", x"71", x"0A", x"A3", x"17", x"D0", x"16",
		x"62", x"14", x"22", x"C1", x"D0", x"16", x"62", x"05", x"22", x"C1", x"75", x"01", x"54", x"50", x"12", x"35",
		x"65", x"00", x"60", x"17", x"61", x"08", x"A3", x"17", x"F3", x"0A", x"33", x"04", x"12", x"79", x"63", x"00",
		x"12", x"97", x"33", x"05", x"12", x"83", x"70", x"0A", x"63", x"01", x"12", x"97", x"33", x"07", x"12", x"8D",
		x"71", x"0A", x"63", x"02", x"12", x"97", x"33", x"08", x"12", x"69", x"70", x"0A", x"71", x"0A", x"63", x"03",
		x"D0", x"16", x"62", x"14", x"22", x"C1", x"D0", x"16", x"A3", x"59", x"F5", x"1E", x"F0", x"65", x"75", x"01",
		x"50", x"30", x"12", x"B5", x"55", x"40", x"12", x"69", x"22", x"DF", x"74", x"01", x"12", x"2D", x"22", x"F9",
		x"A3", x"45", x"60", x"10", x"61", x"0E", x"22", x"CB", x"12", x"BF", x"F2", x"15", x"F2", x"07", x"32", x"00",
		x"12", x"C3", x"00", x"EE", x"83", x"00", x"62", x"05", x"D0", x"15", x"F2", x"1E", x"70", x"08", x"85", x"30",
		x"75", x"20", x"50", x"50", x"12", x"CF", x"00", x"EE", x"A3", x"59", x"83", x"40", x"73", x"FD", x"F3", x"33",
		x"F2", x"65", x"F1", x"29", x"60", x"2B", x"63", x"1B", x"D0", x"35", x"70", x"05", x"F2", x"29", x"D0", x"35",
		x"00", x"EE", x"A3", x"0F", x"60", x"17", x"61", x"07", x"D0", x"18", x"70", x"0A", x"D0", x"18", x"71", x"0A",
		x"D0", x"18", x"70", x"F6", x"D0", x"18", x"00", x"EE", x"FF", x"81", x"81", x"81", x"81", x"81", x"81", x"FF",
		x"7E", x"7E", x"7E", x"7E", x"7E", x"7E", x"DB", x"AA", x"8B", x"CB", x"CB", x"EF", x"08", x"8F", x"0D", x"EC",
		x"A0", x"A0", x"B0", x"30", x"BE", x"5F", x"51", x"51", x"D9", x"D9", x"83", x"82", x"83", x"82", x"FB", x"E8",
		x"08", x"88", x"05", x"E2", x"BE", x"A0", x"B8", x"20", x"3E", x"80", x"80", x"80", x"80", x"F8", x"F7", x"85",
		x"B7", x"95", x"F5", x"76", x"54", x"56", x"54", x"56", x"3A", x"2A", x"2A", x"2A", x"39", x"B6", x"A5", x"B6",
		x"A5", x"35", x"12", x"19", x"4D", x"49", x"53", x"53", x"49", x"4C", x"45", x"20", x"62", x"79", x"20", x"44",
		x"61", x"76", x"69", x"64", x"20", x"57", x"49", x"4E", x"54", x"45", x"52", x"6C", x"0C", x"60", x"00", x"61",
		x"00", x"65", x"08", x"66", x"0A", x"67", x"00", x"6E", x"01", x"A2", x"AD", x"D0", x"14", x"70", x"08", x"30",
		x"40", x"12", x"29", x"60", x"00", x"61", x"1C", x"A2", x"B0", x"D0", x"14", x"A2", x"B0", x"D0", x"14", x"3E",
		x"01", x"12", x"49", x"70", x"04", x"40", x"38", x"6E", x"00", x"12", x"4F", x"70", x"FC", x"40", x"00", x"6E",
		x"01", x"D0", x"14", x"FC", x"15", x"FB", x"07", x"3B", x"00", x"12", x"53", x"62", x"08", x"E2", x"9E", x"12",
		x"95", x"3C", x"00", x"7C", x"FE", x"63", x"1B", x"82", x"00", x"A2", x"B0", x"D2", x"31", x"64", x"00", x"D2",
		x"31", x"73", x"FF", x"D2", x"31", x"3F", x"00", x"64", x"01", x"33", x"03", x"12", x"6D", x"D2", x"31", x"34",
		x"01", x"12", x"91", x"77", x"05", x"75", x"FF", x"82", x"00", x"63", x"00", x"A2", x"AD", x"D2", x"34", x"45",
		x"00", x"12", x"97", x"76", x"FF", x"36", x"00", x"12", x"39", x"A2", x"B4", x"F7", x"33", x"F2", x"65", x"63",
		x"1B", x"64", x"0D", x"F1", x"29", x"D3", x"45", x"73", x"05", x"F2", x"29", x"D3", x"45", x"12", x"AB", x"10",
		x"38", x"38", x"10", x"38", x"7C", x"FE", x"22", x"FC", x"6B", x"0C", x"6C", x"3F", x"6D", x"0C", x"A2", x"EA",
		x"DA", x"B6", x"DC", x"D6", x"6E", x"00", x"22", x"D4", x"66", x"03", x"68", x"02", x"60", x"60", x"F0", x"15",
		x"F0", x"07", x"30", x"00", x"12", x"1A", x"C7", x"17", x"77", x"08", x"69", x"FF", x"A2", x"F0", x"D6", x"71",
		x"A2", x"EA", x"DA", x"B6", x"DC", x"D6", x"60", x"01", x"E0", x"A1", x"7B", x"FE", x"60", x"04", x"E0", x"A1",
		x"7B", x"02", x"60", x"1F", x"8B", x"02", x"DA", x"B6", x"60", x"0C", x"E0", x"A1", x"7D", x"FE", x"60", x"0D",
		x"E0", x"A1", x"7D", x"02", x"60", x"1F", x"8D", x"02", x"DC", x"D6", x"A2", x"F0", x"D6", x"71", x"86", x"84",
		x"87", x"94", x"60", x"3F", x"86", x"02", x"61", x"1F", x"87", x"12", x"46", x"00", x"12", x"78", x"46", x"3F",
		x"12", x"82", x"47", x"1F", x"69", x"FF", x"47", x"00", x"69", x"01", x"D6", x"71", x"12", x"2A", x"68", x"02",
		x"63", x"01", x"80", x"70", x"80", x"B5", x"12", x"8A", x"68", x"FE", x"63", x"0A", x"80", x"70", x"80", x"D5",
		x"3F", x"01", x"12", x"A2", x"61", x"02", x"80", x"15", x"3F", x"01", x"12", x"BA", x"80", x"15", x"3F", x"01",
		x"12", x"C8", x"80", x"15", x"3F", x"01", x"12", x"C2", x"60", x"20", x"F0", x"18", x"22", x"D4", x"8E", x"34",
		x"22", x"D4", x"66", x"3E", x"33", x"01", x"66", x"03", x"68", x"FE", x"33", x"01", x"68", x"02", x"12", x"16",
		x"79", x"FF", x"49", x"FE", x"69", x"FF", x"12", x"C8", x"79", x"01", x"49", x"02", x"69", x"01", x"60", x"04",
		x"F0", x"18", x"76", x"01", x"46", x"40", x"76", x"FE", x"12", x"6C", x"A2", x"F2", x"FE", x"33", x"F2", x"65",
		x"F1", x"29", x"64", x"14", x"65", x"02", x"D4", x"55", x"74", x"15", x"F2", x"29", x"D4", x"55", x"00", x"EE",
		x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00", x"00", x"00", x"C0", x"C0", x"C0", x"00",
		x"FF", x"00", x"6B", x"20", x"6C", x"00", x"A2", x"F6", x"DB", x"C4", x"7C", x"04", x"3C", x"20", x"13", x"02",
		x"6A", x"00", x"6B", x"00", x"6C", x"1F", x"A2", x"FA", x"DA", x"B1", x"DA", x"C1", x"7A", x"08", x"3A", x"40",
		x"13", x"12", x"A2", x"F6", x"6A", x"00", x"6B", x"20", x"DB", x"A1", x"00", x"EE", x"22", x"F6", x"6B", x"0C",
		x"6C", x"3F", x"6D", x"0C", x"A2", x"EA", x"DA", x"B6", x"DC", x"D6", x"6E", x"00", x"22", x"D4", x"66", x"03",
		x"68", x"02", x"60", x"60", x"F0", x"15", x"F0", x"07", x"30", x"00", x"12", x"1A", x"C7", x"17", x"77", x"08",
		x"69", x"FF", x"A2", x"F0", x"D6", x"71", x"A2", x"EA", x"DA", x"B6", x"DC", x"D6", x"60", x"01", x"E0", x"A1",
		x"7B", x"FE", x"60", x"04", x"E0", x"A1", x"7B", x"02", x"60", x"1F", x"8B", x"02", x"DA", x"B6", x"60", x"0C",
		x"E0", x"A1", x"7D", x"FE", x"60", x"0D", x"E0", x"A1", x"7D", x"02", x"60", x"1F", x"8D", x"02", x"DC", x"D6",
		x"A2", x"F0", x"D6", x"71", x"86", x"84", x"87", x"94", x"60", x"3F", x"86", x"02", x"61", x"1F", x"87", x"12",
		x"46", x"00", x"12", x"78", x"46", x"3F", x"12", x"82", x"47", x"1F", x"69", x"FF", x"47", x"00", x"69", x"01",
		x"D6", x"71", x"12", x"2A", x"68", x"02", x"63", x"01", x"80", x"70", x"80", x"B5", x"12", x"8A", x"68", x"FE",
		x"63", x"0A", x"80", x"70", x"80", x"D5", x"3F", x"01", x"12", x"A2", x"61", x"02", x"80", x"15", x"3F", x"01",
		x"12", x"BA", x"80", x"15", x"3F", x"01", x"12", x"C8", x"80", x"15", x"3F", x"01", x"12", x"C2", x"60", x"20",
		x"F0", x"18", x"22", x"D4", x"8E", x"34", x"22", x"D4", x"66", x"3E", x"33", x"01", x"66", x"03", x"68", x"FE",
		x"33", x"01", x"68", x"02", x"12", x"16", x"79", x"FF", x"49", x"FE", x"69", x"FF", x"12", x"C8", x"79", x"01",
		x"49", x"02", x"69", x"01", x"60", x"04", x"F0", x"18", x"76", x"01", x"46", x"40", x"76", x"FE", x"12", x"6C",
		x"A2", x"F2", x"FE", x"33", x"F2", x"65", x"F1", x"29", x"64", x"14", x"65", x"00", x"D4", x"55", x"74", x"15",
		x"F2", x"29", x"D4", x"55", x"00", x"EE", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"00", x"00", x"00",
		x"00", x"00", x"6B", x"20", x"6C", x"00", x"A2", x"EA", x"DB", x"C1", x"7C", x"01", x"3C", x"20", x"12", x"FC",
		x"6A", x"00", x"00", x"EE", x"6A", x"12", x"6B", x"01", x"61", x"10", x"62", x"00", x"60", x"00", x"A2", x"B0",
		x"D1", x"27", x"F0", x"29", x"30", x"00", x"DA", x"B5", x"71", x"08", x"7A", x"08", x"31", x"30", x"12", x"24",
		x"61", x"10", x"72", x"08", x"6A", x"12", x"7B", x"08", x"A3", x"00", x"F0", x"1E", x"F0", x"55", x"70", x"01",
		x"30", x"10", x"12", x"0A", x"6A", x"12", x"6B", x"01", x"6C", x"00", x"62", x"FF", x"C0", x"06", x"70", x"02",
		x"22", x"52", x"72", x"FF", x"32", x"00", x"12", x"38", x"6E", x"00", x"6E", x"00", x"F0", x"0A", x"22", x"52",
		x"7E", x"01", x"7E", x"01", x"12", x"48", x"84", x"A0", x"85", x"B0", x"86", x"C0", x"30", x"02", x"12", x"64",
		x"45", x"01", x"12", x"64", x"75", x"F8", x"76", x"FC", x"30", x"08", x"12", x"70", x"45", x"19", x"12", x"70",
		x"75", x"08", x"76", x"04", x"30", x"06", x"12", x"7C", x"44", x"12", x"12", x"7C", x"74", x"F8", x"76", x"FF",
		x"30", x"04", x"12", x"88", x"44", x"2A", x"12", x"88", x"74", x"08", x"76", x"01", x"A3", x"00", x"F6", x"1E",
		x"F0", x"65", x"81", x"00", x"60", x"00", x"A3", x"00", x"F6", x"1E", x"F0", x"55", x"A3", x"00", x"FC", x"1E",
		x"80", x"10", x"F0", x"55", x"F1", x"29", x"D4", x"55", x"DA", x"B5", x"8A", x"40", x"8B", x"50", x"8C", x"60",
		x"00", x"EE", x"EE", x"5E", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"FE", x"6D", x"02", x"6E", x"02",
		x"6C", x"00", x"A2", x"D7", x"6B", x"00", x"6A", x"11", x"DA", x"B3", x"3A", x"2D", x"12", x"1A", x"4B", x"1C",
		x"12", x"1E", x"7B", x"04", x"12", x"0A", x"7A", x"04", x"12", x"0C", x"6A", x"1D", x"6B", x"0C", x"DA", x"B3",
		x"7A", x"04", x"7B", x"04", x"DA", x"B3", x"A2", x"DA", x"DA", x"B3", x"7A", x"FC", x"DA", x"B3", x"7B", x"FC",
		x"DA", x"B3", x"7A", x"04", x"DA", x"B3", x"60", x"02", x"22", x"DE", x"60", x"34", x"22", x"DE", x"A2", x"D7",
		x"60", x"34", x"22", x"DE", x"23", x"94", x"69", x"01", x"23", x"0C", x"68", x"00", x"23", x"7E", x"69", x"00",
		x"49", x"09", x"12", x"72", x"79", x"01", x"E9", x"9E", x"12", x"54", x"49", x"05", x"12", x"8C", x"38", x"00",
		x"23", x"9E", x"23", x"0C", x"38", x"00", x"23", x"9E", x"61", x"02", x"F1", x"18", x"12", x"50", x"69", x"0F",
		x"E9", x"9E", x"12", x"50", x"38", x"00", x"22", x"EC", x"7C", x"80", x"38", x"00", x"22", x"EC", x"61", x"18",
		x"F1", x"18", x"E9", x"A1", x"12", x"86", x"12", x"50", x"38", x"00", x"23", x"7E", x"23", x"A8", x"31", x"00",
		x"12", x"50", x"83", x"A0", x"84", x"B0", x"69", x"00", x"23", x"D0", x"42", x"00", x"12", x"50", x"23", x"94",
		x"A2", x"DA", x"D3", x"43", x"3C", x"00", x"12", x"B0", x"A2", x"D7", x"D3", x"43", x"3C", x"00", x"12", x"B8",
		x"7D", x"01", x"12", x"BA", x"7E", x"01", x"23", x"FA", x"23", x"D0", x"32", x"00", x"12", x"BA", x"23", x"94",
		x"81", x"D0", x"81", x"E4", x"31", x"40", x"12", x"78", x"24", x"2E", x"24", x"2E", x"23", x"88", x"24", x"2E",
		x"12", x"CC", x"01", x"00", x"40", x"00", x"E0", x"A0", x"E0", x"D4", x"61", x"0B", x"D0", x"13", x"70", x"04",
		x"D0", x"73", x"70", x"04", x"D0", x"13", x"00", x"EE", x"A4", x"40", x"3C", x"00", x"13", x"06", x"65", x"02",
		x"FD", x"33", x"66", x"04", x"F2", x"65", x"F1", x"29", x"D5", x"65", x"75", x"07", x"F2", x"29", x"D5", x"65",
		x"00", x"EE", x"65", x"34", x"FE", x"33", x"12", x"F6", x"67", x"00", x"49", x"09", x"13", x"72", x"49", x"08",
		x"13", x"5E", x"49", x"07", x"13", x"66", x"49", x"06", x"13", x"56", x"49", x"04", x"13", x"4E", x"49", x"03",
		x"13", x"42", x"49", x"01", x"13", x"36", x"4B", x"00", x"13", x"32", x"7B", x"FC", x"00", x"EE", x"67", x"FF",
		x"00", x"EE", x"4B", x"00", x"13", x"32", x"4A", x"11", x"13", x"32", x"7A", x"FC", x"13", x"2E", x"4B", x"00",
		x"13", x"32", x"4A", x"2D", x"13", x"32", x"7A", x"04", x"13", x"2E", x"4A", x"11", x"13", x"32", x"7A", x"FC",
		x"00", x"EE", x"4A", x"2D", x"13", x"32", x"7A", x"04", x"00", x"EE", x"4B", x"1C", x"13", x"32", x"7B", x"04",
		x"00", x"EE", x"4B", x"1C", x"13", x"32", x"4A", x"11", x"13", x"32", x"7A", x"FC", x"13", x"62", x"4B", x"1C",
		x"13", x"32", x"4A", x"2D", x"13", x"32", x"7A", x"04", x"13", x"62", x"23", x"88", x"22", x"EC", x"23", x"9E",
		x"78", x"80", x"00", x"EE", x"61", x"10", x"F1", x"15", x"F1", x"07", x"31", x"00", x"13", x"8C", x"00", x"EE",
		x"22", x"EC", x"7C", x"80", x"22", x"EC", x"7C", x"80", x"00", x"EE", x"A2", x"D7", x"DA", x"B3", x"00", x"EE",
		x"A2", x"DA", x"13", x"A0", x"23", x"A4", x"81", x"F0", x"23", x"A4", x"41", x"00", x"13", x"CC", x"23", x"9E",
		x"81", x"F0", x"23", x"9E", x"31", x"00", x"13", x"C4", x"3C", x"00", x"13", x"C8", x"61", x"80", x"00", x"EE",
		x"3C", x"00", x"13", x"C0", x"61", x"FF", x"00", x"EE", x"61", x"00", x"00", x"EE", x"8A", x"30", x"8B", x"40",
		x"79", x"01", x"49", x"05", x"79", x"01", x"62", x"00", x"49", x"0A", x"00", x"EE", x"23", x"0C", x"23", x"A8",
		x"41", x"00", x"13", x"D0", x"31", x"80", x"13", x"F2", x"32", x"00", x"00", x"EE", x"13", x"D0", x"47", x"FF",
		x"13", x"D0", x"72", x"01", x"13", x"E0", x"81", x"90", x"69", x"0A", x"89", x"15", x"23", x"0C", x"81", x"A0",
		x"81", x"35", x"31", x"00", x"14", x"1A", x"81", x"B0", x"81", x"45", x"31", x"00", x"14", x"1A", x"81", x"90",
		x"69", x"0A", x"89", x"15", x"00", x"EE", x"23", x"9E", x"3C", x"00", x"14", x"26", x"7D", x"01", x"7E", x"FF",
		x"14", x"2A", x"7D", x"FF", x"7E", x"01", x"24", x"2E", x"14", x"00", x"61", x"04", x"F1", x"18", x"23", x"88",
		x"00", x"EE", x"14", x"24", x"4A", x"2D", x"14", x"24", x"7A", x"04", x"14", x"20", x"00", x"00", x"00", x"E0",
		x"C0", x"FF", x"A2", x"24", x"F0", x"33", x"F2", x"65", x"F0", x"29", x"60", x"00", x"63", x"00", x"D0", x"35",
		x"F1", x"29", x"60", x"05", x"D0", x"35", x"F2", x"29", x"60", x"0A", x"D0", x"35", x"F0", x"0A", x"12", x"00",
		x"2D", x"47", x"50", x"10", x"2F", x"0E", x"12", x"24", x"5B", x"62", x"79", x"20", x"68", x"61", x"70", x"5D",
		x"9A", x"00", x"88", x"00", x"84", x"35", x"88", x"00", x"88", x"6A", x"80", x"27", x"84", x"35", x"80", x"27",
		x"88", x"6A", x"84", x"19", x"00", x"E0", x"A8", x"96", x"FA", x"65", x"F3", x"15", x"A8", x"97", x"F2", x"1E",
		x"F1", x"65", x"A8", x"75", x"F0", x"1E", x"24", x"B3", x"D4", x"A7", x"F1", x"1E", x"D9", x"A7", x"FA", x"18",
		x"74", x"08", x"79", x"F8", x"72", x"02", x"32", x"08", x"12", x"2A", x"60", x"0A", x"24", x"B1", x"68", x"48",
		x"2D", x"BD", x"2D", x"47", x"50", x"10", x"1F", x"2C", x"24", x"AF", x"68", x"5D", x"2D", x"BD", x"F0", x"0A",
		x"00", x"E0", x"60", x"0F", x"24", x"B1", x"A8", x"92", x"F1", x"65", x"A4", x"25", x"F1", x"55", x"A7", x"F7",
		x"F5", x"65", x"A8", x"29", x"D5", x"46", x"75", x"08", x"35", x"40", x"12", x"74", x"D4", x"0D", x"D4", x"1C",
		x"74", x"08", x"34", x"28", x"12", x"7C", x"72", x"06", x"61", x"08", x"A7", x"9A", x"42", x"20", x"A7", x"96",
		x"D2", x"15", x"A8", x"03", x"F3", x"1E", x"73", x"01", x"F0", x"65", x"A7", x"FC", x"30", x"00", x"D2", x"14",
		x"42", x"20", x"12", x"C2", x"61", x"07", x"A8", x"03", x"F3", x"1E", x"F0", x"65", x"71", x"06", x"41", x"1F",
		x"12", x"86", x"A7", x"95", x"D2", x"16", x"40", x"00", x"12", x"AC", x"A7", x"FB", x"D2", x"15", x"70", x"FF",
		x"12", x"AC", x"68", x"36", x"2D", x"BD", x"A8", x"89", x"FE", x"65", x"67", x"0A", x"23", x"41", x"A7", x"8F",
		x"D7", x"B1", x"24", x"B3", x"F9", x"0A", x"D7", x"B1", x"49", x"01", x"13", x"8B", x"49", x"0A", x"13", x"99",
		x"60", x"06", x"F0", x"15", x"23", x"49", x"66", x"00", x"49", x"05", x"13", x"06", x"49", x"08", x"13", x"14",
		x"49", x"09", x"13", x"24", x"39", x"07", x"12", x"CC", x"47", x"0A", x"12", x"CC", x"7C", x"FF", x"77", x"FA",
		x"66", x"FF", x"65", x"74", x"13", x"36", x"4B", x"0A", x"12", x"CC", x"7D", x"FF", x"7B", x"FA", x"66", x"FF",
		x"65", x"BA", x"13", x"38", x"4B", x"1C", x"12", x"CC", x"47", x"22", x"12", x"CC", x"7D", x"01", x"7B", x"06",
		x"65", x"46", x"13", x"38", x"47", x"22", x"12", x"CC", x"37", x"1C", x"13", x"30", x"3B", x"0A", x"12", x"CC",
		x"7C", x"01", x"77", x"06", x"65", x"8C", x"23", x"6F", x"23", x"6F", x"12", x"CC", x"36", x"3B", x"08", x"2C",
		x"31", x"80", x"C0", x"81", x"D0", x"A7", x"ED", x"F1", x"55", x"A3", x"3C", x"F4", x"65", x"4E", x"00", x"13",
		x"61", x"A2", x"61", x"D0", x"21", x"72", x"FE", x"80", x"E0", x"40", x"0A", x"60", x"0F", x"F0", x"29", x"D1",
		x"25", x"A7", x"ED", x"F1", x"65", x"F1", x"29", x"D4", x"25", x"F0", x"29", x"D3", x"25", x"00", x"EE", x"A4",
		x"25", x"F1", x"65", x"82", x"60", x"81", x"54", x"4F", x"01", x"13", x"81", x"46", x"FF", x"70", x"FF", x"13",
		x"85", x"46", x"00", x"70", x"01", x"A4", x"25", x"F1", x"55", x"00", x"EE", x"2D", x"55", x"F9", x"18", x"68",
		x"2F", x"2D", x"BD", x"60", x"2D", x"24", x"B1", x"12", x"24", x"4F", x"01", x"13", x"B1", x"2D", x"55", x"F9",
		x"18", x"68", x"28", x"2D", x"BD", x"60", x"2D", x"24", x"B1", x"68", x"28", x"2D", x"BD", x"2D", x"55", x"12",
		x"CE", x"2D", x"55", x"24", x"A7", x"7E", x"01", x"00", x"E0", x"2D", x"55", x"68", x"00", x"2D", x"BD", x"23",
		x"49", x"88", x"E0", x"78", x"FF", x"80", x"0E", x"88", x"04", x"88", x"22", x"88", x"8E", x"A2", x"0C", x"F7",
		x"65", x"A2", x"14", x"F8", x"1E", x"F3", x"65", x"85", x"10", x"87", x"30", x"A2", x"0C", x"F7", x"55", x"A7",
		x"E0", x"FC", x"65", x"A6", x"9C", x"F1", x"55", x"A6", x"A2", x"F1", x"55", x"A8", x"58", x"24", x"6B", x"62",
		x"0F", x"A8", x"69", x"24", x"6B", x"FC", x"29", x"D3", x"55", x"73", x"05", x"33", x"40", x"13", x"F7", x"A7",
		x"AC", x"D4", x"CA", x"D4", x"6A", x"D4", x"5C", x"DC", x"CA", x"DC", x"6A", x"DC", x"5C", x"A8", x"29", x"D7",
		x"AF", x"D7", x"8F", x"77", x"08", x"37", x"24", x"14", x"0F", x"A7", x"8E", x"D4", x"67", x"68", x"FF", x"3B",
		x"00", x"14", x"2F", x"6B", x"08", x"A8", x"A1", x"FC", x"1E", x"F0", x"65", x"8D", x"00", x"7C", x"01", x"7B",
		x"FF", x"8D", x"D6", x"4F", x"00", x"14", x"3D", x"78", x"01", x"38", x"03", x"14", x"1F", x"48", x"FF", x"14",
		x"55", x"4A", x"0B", x"78", x"04", x"24", x"7D", x"88", x"86", x"4F", x"01", x"14", x"55", x"79", x"FD", x"88",
		x"86", x"4F", x"01", x"79", x"05", x"79", x"05", x"39", x"23", x"14", x"1D", x"69", x"05", x"7A", x"05", x"3A",
		x"1F", x"14", x"1D", x"A7", x"E4", x"FD", x"65", x"2D", x"BD", x"14", x"E7", x"60", x"29", x"D0", x"24", x"70",
		x"08", x"40", x"41", x"00", x"EE", x"F7", x"1E", x"14", x"6D", x"2D", x"1F", x"1B", x"24", x"A2", x"0B", x"F8",
		x"1E", x"F1", x"65", x"80", x"80", x"80", x"06", x"4F", x"01", x"14", x"9F", x"A4", x"79", x"F0", x"1E", x"F0",
		x"65", x"A7", x"9E", x"F1", x"1E", x"D9", x"A5", x"F0", x"1E", x"79", x"08", x"D9", x"A5", x"00", x"EE", x"A7",
		x"9E", x"F1", x"1E", x"D9", x"AF", x"00", x"EE", x"60", x"01", x"F0", x"18", x"68", x"23", x"2D", x"BD", x"60",
		x"21", x"F0", x"15", x"F0", x"07", x"30", x"00", x"14", x"B3", x"00", x"EE", x"E5", x"A1", x"14", x"BB", x"A7",
		x"FF", x"DB", x"C5", x"2D", x"55", x"68", x"12", x"2D", x"BD", x"F9", x"0A", x"68", x"12", x"2D", x"BD", x"39",
		x"0A", x"14", x"D7", x"24", x"A7", x"13", x"B7", x"2D", x"BD", x"F9", x"0A", x"68", x"1B", x"2D", x"BD", x"39",
		x"0A", x"14", x"E7", x"24", x"A7", x"12", x"60", x"2D", x"55", x"15", x"41", x"25", x"C5", x"15", x"41", x"25",
		x"97", x"26", x"21", x"14", x"FF", x"25", x"F1", x"25", x"97", x"15", x"41", x"25", x"C5", x"26", x"21", x"3B",
		x"FF", x"15", x"41", x"66", x"00", x"65", x"07", x"23", x"6F", x"3E", x"0A", x"13", x"B5", x"00", x"E0", x"68",
		x"6B", x"2D", x"BD", x"A7", x"EC", x"F2", x"65", x"41", x"05", x"15", x"3B", x"A8", x"03", x"F1", x"1E", x"F0",
		x"65", x"40", x"03", x"15", x"3B", x"72", x"F6", x"50", x"20", x"15", x"3B", x"70", x"01", x"A8", x"03", x"F1",
		x"1E", x"F0", x"55", x"2D", x"BD", x"2D", x"47", x"50", x"10", x"2E", x"CE", x"12", x"58", x"25", x"C5", x"25",
		x"F1", x"A7", x"FF", x"DB", x"C5", x"A7", x"F1", x"F6", x"65", x"E5", x"A1", x"14", x"BB", x"E2", x"A1", x"70",
		x"02", x"E1", x"A1", x"70", x"04", x"E3", x"A1", x"70", x"08", x"E6", x"A1", x"70", x"10", x"40", x"00", x"15",
		x"93", x"FA", x"07", x"3A", x"00", x"15", x"45", x"F4", x"15", x"E4", x"A1", x"65", x"02", x"A7", x"FF", x"DB",
		x"C5", x"85", x"F1", x"B5", x"73", x"14", x"F7", x"14", x"FD", x"14", x"EF", x"14", x"EB", x"14", x"F7", x"14",
		x"FB", x"14", x"EF", x"15", x"3F", x"14", x"F5", x"14", x"FD", x"14", x"EF", x"15", x"3D", x"14", x"F5", x"14",
		x"FB", x"14", x"EF", x"F0", x"15", x"15", x"45", x"4B", x"23", x"00", x"EE", x"4C", x"01", x"00", x"EE", x"35",
		x"03", x"15", x"C1", x"27", x"02", x"9A", x"90", x"00", x"EE", x"80", x"A0", x"70", x"FF", x"A8", x"17", x"DB",
		x"01", x"DB", x"01", x"4F", x"01", x"00", x"EE", x"89", x"B0", x"24", x"7D", x"7A", x"FB", x"24", x"7D", x"26",
		x"A6", x"7C", x"FB", x"00", x"EE", x"4B", x"23", x"00", x"EE", x"4C", x"1A", x"00", x"EE", x"35", x"03", x"15",
		x"ED", x"27", x"02", x"9A", x"90", x"00", x"EE", x"79", x"05", x"A8", x"17", x"DB", x"91", x"DB", x"91", x"4F",
		x"01", x"00", x"EE", x"89", x"B0", x"24", x"7D", x"7A", x"05", x"24", x"7D", x"26", x"A6", x"7C", x"05", x"00",
		x"EE", x"4B", x"05", x"00", x"EE", x"35", x"03", x"16", x"17", x"27", x"46", x"99", x"60", x"00", x"EE", x"80",
		x"90", x"70", x"FF", x"A8", x"18", x"D0", x"C3", x"D0", x"C3", x"4F", x"01", x"00", x"EE", x"8A", x"C0", x"24",
		x"7D", x"79", x"F3", x"24", x"7D", x"26", x"A6", x"7B", x"FB", x"00", x"EE", x"4C", x"0B", x"16", x"29", x"00",
		x"EE", x"4B", x"1E", x"16", x"1B", x"4B", x"23", x"00", x"EE", x"35", x"03", x"16", x"4D", x"27", x"46", x"99",
		x"60", x"00", x"EE", x"76", x"05", x"A8", x"18", x"D6", x"C3", x"D6", x"C3", x"4F", x"01", x"00", x"EE", x"8A",
		x"C0", x"24", x"7D", x"79", x"FD", x"24", x"7D", x"26", x"A6", x"46", x"23", x"16", x"51", x"7B", x"05", x"00",
		x"EE", x"7B", x"05", x"86", x"B0", x"8B", x"90", x"7B", x"F3", x"A8", x"17", x"DB", x"C1", x"DB", x"C1", x"4F",
		x"00", x"16", x"6D", x"A8", x"13", x"DB", x"C5", x"DB", x"C5", x"4F", x"01", x"16", x"83", x"4B", x"05", x"16",
		x"75", x"7B", x"FB", x"16", x"59", x"87", x"80", x"2D", x"55", x"68", x"0A", x"2D", x"BD", x"6A", x"0B", x"88",
		x"70", x"66", x"FF", x"63", x"00", x"8B", x"60", x"62", x"0B", x"F2", x"18", x"F2", x"15", x"79", x"F8", x"24",
		x"7D", x"73", x"01", x"24", x"B3", x"33", x"0B", x"16", x"8B", x"00", x"EE", x"00", x"00", x"00", x"36", x"3B",
		x"14", x"00", x"00", x"00", x"2C", x"31", x"A6", x"9C", x"F4", x"65", x"F5", x"18", x"7D", x"01", x"A6", x"9B",
		x"FD", x"33", x"41", x"09", x"16", x"C2", x"F1", x"29", x"D3", x"45", x"71", x"01", x"F1", x"29", x"D3", x"45",
		x"00", x"EE", x"F0", x"29", x"D2", x"45", x"F1", x"29", x"D3", x"45", x"A6", x"9C", x"F1", x"65", x"F0", x"29",
		x"D2", x"45", x"F1", x"29", x"D3", x"45", x"4D", x"64", x"16", x"DC", x"00", x"EE", x"A6", x"A2", x"F3", x"65",
		x"6D", x"00", x"77", x"01", x"47", x"64", x"67", x"00", x"A6", x"A1", x"F7", x"33", x"F0", x"29", x"D2", x"45",
		x"F1", x"29", x"D3", x"45", x"A6", x"A2", x"F1", x"65", x"F0", x"29", x"D2", x"45", x"F1", x"29", x"D3", x"45",
		x"00", x"EE", x"68", x"01", x"8A", x"C0", x"89", x"C0", x"A8", x"13", x"DB", x"95", x"DB", x"95", x"4F", x"01",
		x"17", x"22", x"79", x"05", x"DB", x"95", x"DB", x"95", x"4F", x"01", x"17", x"22", x"79", x"05", x"78", x"02",
		x"00", x"EE", x"A8", x"17", x"DB", x"A1", x"DB", x"A1", x"4F", x"01", x"17", x"3C", x"7A", x"FB", x"DB", x"A1",
		x"DB", x"A1", x"4F", x"01", x"17", x"3C", x"7A", x"FB", x"78", x"02", x"00", x"EE", x"80", x"90", x"80", x"A5",
		x"40", x"0A", x"78", x"02", x"00", x"EE", x"68", x"00", x"4C", x"0B", x"78", x"04", x"89", x"B0", x"86", x"B0",
		x"A8", x"1B", x"D6", x"C3", x"D6", x"C3", x"4F", x"01", x"17", x"6A", x"76", x"05", x"D6", x"C3", x"D6", x"C3",
		x"4F", x"01", x"17", x"6A", x"76", x"05", x"78", x"02", x"00", x"EE", x"A8", x"18", x"D9", x"C3", x"D9", x"C3",
		x"4F", x"01", x"17", x"84", x"79", x"FB", x"D9", x"C3", x"D9", x"C3", x"4F", x"01", x"17", x"84", x"79", x"FB",
		x"78", x"02", x"00", x"EE", x"80", x"60", x"80", x"95", x"40", x"0A", x"78", x"02", x"00", x"EE", x"D0", x"80",
		x"80", x"80", x"80", x"80", x"D0", x"20", x"F8", x"88", x"88", x"88", x"F8", x"88", x"8C", x"88", x"F8", x"D8",
		x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"F8", x"F8", x"F8", x"F8",
		x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"F8", x"88", x"A8", x"A8", x"88", x"88", x"A8", x"A8", x"A8",
		x"88", x"88", x"A8", x"A8", x"88", x"F8", x"88", x"C8", x"A8", x"98", x"88", x"C8", x"A8", x"98", x"88", x"C8",
		x"A8", x"98", x"88", x"F8", x"88", x"A8", x"A8", x"88", x"88", x"A8", x"A8", x"88", x"F8", x"00", x"00", x"00",
		x"00", x"00", x"01", x"2C", x"23", x"14", x"0A", x"04", x"10", x"05", x"01", x"00", x"00", x"00", x"00", x"05",
		x"01", x"00", x"09", x"05", x"08", x"0A", x"01", x"07", x"14", x"02", x"00", x"00", x"00", x"70", x"70", x"70",
		x"F8", x"F8", x"F8", x"70", x"00", x"00", x"00", x"00", x"F8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8", x"D8",
		x"D8", x"F8", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"00", x"80", x"00", x"00", x"08", x"FF", x"88",
		x"91", x"A2", x"FF", x"80", x"B3", x"80", x"FF", x"FF", x"80", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF",
		x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FD", x"FC", x"80", x"FC", x"FD", x"FE", x"8A", x"12",
		x"22", x"FE", x"02", x"9A", x"02", x"FE", x"FE", x"02", x"FE", x"FE", x"EE", x"E6", x"02", x"E6", x"EE", x"C0",
		x"40", x"40", x"40", x"C0", x"C0", x"40", x"C0", x"C0", x"83", x"E4", x"94", x"E3", x"33", x"8A", x"AA", x"1A",
		x"08", x"38", x"48", x"38", x"38", x"38", x"38", x"38", x"38", x"F1", x"AA", x"AA", x"A9", x"94", x"55", x"49",
		x"88", x"8C", x"50", x"04", x"D8", x"FC", x"E6", x"E6", x"E4", x"F8", x"EC", x"E6", x"E6", x"E6", x"FE", x"E6",
		x"E6", x"E6", x"E6", x"E6", x"E6", x"7C", x"E6", x"E0", x"7C", x"06", x"E6", x"7C", x"E6", x"E6", x"E6", x"E6",
		x"E6", x"7C", x"A8", x"A1", x"0A", x"01", x"0A", x"00", x"00", x"0A", x"00", x"10", x"06", x"06", x"00", x"39",
		x"01", x"E1", x"9F", x"47", x"00", x"86", x"38", x"00", x"E3", x"30", x"1F", x"73", x"60", x"4A", x"00", x"00",
		x"A0", x"47", x"BC", x"01", x"01", x"00", x"CF", x"03", x"08", x"EC", x"C0", x"38", x"00", x"79", x"7B", x"3C",
		x"31", x"C7", x"10", x"04", x"19", x"F1", x"AF", x"A7", x"61", x"00", x"07", x"D6", x"86", x"21", x"46", x"60",
		x"00", x"00", x"E8", x"69", x"DA", x"88", x"DA", x"E5", x"00", x"56", x"58", x"F1", x"FB", x"83", x"31", x"00",
		x"4D", x"E1", x"3F", x"38", x"B0", x"22", x"00", x"DF", x"03", x"08", x"EC", x"C0", x"38", x"00", x"8B", x"E7",
		x"11", x"E0", x"60", x"0E", x"00", x"35", x"8C", x"37", x"79", x"82", x"25", x"01", x"0D", x"D0", x"D6", x"46",
		x"30", x"05", x"00", x"4A", x"FD", x"FF", x"07", x"1B", x"90", x"02", x"B5", x"9F", x"B0", x"0F", x"0E", x"08",
		x"00", x"3B", x"A8", x"86", x"3C", x"67", x"3B", x"00", x"ED", x"09", x"3E", x"38", x"84", x"03", x"00", x"2C",
		x"30", x"16", x"34", x"0E", x"00", x"00", x"E3", x"34", x"1A", x"0F", x"B0", x"E0", x"00", x"ED", x"79", x"20",
		x"38", x"00", x"1C", x"00", x"EC", x"C6", x"27", x"18", x"4D", x"E6", x"00", x"DC", x"B3", x"20", x"6C", x"41",
		x"1C", x"00", x"2C", x"06", x"D3", x"08", x"67", x"02", x"00", x"4D", x"E1", x"3F", x"E3", x"30", x"0B", x"02",
		x"E6", x"C6", x"9E", x"D8", x"0E", x"C6", x"10", x"EB", x"11", x"1A", x"8F", x"30", x"E0", x"00", x"37", x"78",
		x"05", x"9B", x"9E", x"53", x"00", x"E7", x"31", x"84", x"AD", x"68", x"76", x"00", x"6F", x"87", x"21", x"94",
		x"07", x"0A", x"00", x"39", x"AC", x"C5", x"F3", x"09", x"70", x"00", x"FD", x"02", x"82", x"D5", x"63", x"04",
		x"00", x"F6", x"02", x"82", x"D5", x"6B", x"73", x"00", x"E3", x"30", x"1F", x"73", x"83", x"29", x"01", x"7C",
		x"8F", x"11", x"EC", x"D0", x"26", x"00", x"7F", x"59", x"9E", x"B8", x"C1", x"14", x"00", x"4D", x"F1", x"FF",
		x"C1", x"81", x"15", x"01", x"E3", x"34", x"1A", x"8F", x"B0", x"E0", x"00", x"EC", x"30", x"1A", x"9F", x"6C",
		x"41", x"00", x"9F", x"B1", x"F1", x"C8", x"0D", x"A6", x"04", x"7A", x"C0", x"2F", x"F0", x"01", x"10", x"00",
		x"EC", x"F0", x"09", x"46", x"93", x"39", x"00", x"0D", x"A6", x"7F", x"61", x"C1", x"56", x"00", x"F7", x"1B",
		x"43", x"4C", x"D9", x"08", x"0E", x"E6", x"9E", x"8D", x"A0", x"9E", x"25", x"00", x"EC", x"62", x"16", x"6C",
		x"3D", x"E2", x"00", x"67", x"DB", x"C1", x"B7", x"00", x"EB", x"00", x"EA", x"0F", x"2C", x"59", x"07", x"0A",
		x"00", x"DE", x"1A", x"36", x"62", x"CD", x"18", x"70", x"5A", x"62", x"7C", x"C2", x"0F", x"28", x"00", x"6D",
		x"0C", x"69", x"D3", x"80", x"D6", x"01", x"F6", x"82", x"D2", x"EF", x"D0", x"80", x"00", x"EB", x"07", x"68",
		x"30", x"C7", x"5A", x"00", x"73", x"03", x"FA", x"6D", x"C1", x"E6", x"28", x"BB", x"E7", x"68", x"03", x"E2",
		x"86", x"00", x"BF", x"F5", x"30", x"1A", x"4C", x"18", x"07", x"0D", x"3F", x"FE", x"09", x"07", x"56", x"04",
		x"DF", x"C6", x"F0", x"C8", x"0D", x"A6", x"04", x"4B", x"EA", x"63", x"2C", x"D8", x"0A", x"00", x"D6", x"30",
		x"16", x"B4", x"7E", x"84", x"03", x"6B", x"DE", x"80", x"A6", x"1F", x"50", x"02", x"D3", x"73", x"B4", x"01",
		x"71", x"E3", x"00", x"56", x"64", x"6D", x"40", x"D3", x"E6", x"00", x"6B", x"81", x"B5", x"64", x"2D", x"E0",
		x"00", x"2B", x"EC", x"F2", x"B6", x"8C", x"61", x"1C", x"BF", x"1B", x"3C", x"B1", x"06", x"1C", x"05", x"B7",
		x"11", x"BE", x"C1", x"84", x"76", x"00", x"6A", x"6C", x"84", x"7F", x"0B", x"A2", x"03", x"3B", x"D8", x"17",
		x"D6", x"60", x"18", x"07", x"5B", x"1E", x"E8", x"93", x"35", x"8C", x"03", x"5B", x"F1", x"4A", x"9F", x"B1",
		x"80", x"03", x"56", x"AC", x"0F", x"BE", x"01", x"39", x"00", x"F3", x"82", x"7D", x"60", x"67", x"2C", x"01",
		x"2E", x"D6", x"92", x"B5", x"BD", x"D0", x"01", x"B7", x"2D", x"C8", x"58", x"62", x"2D", x"00", x"0A", x"3F",
		x"82", x"AC", x"C5", x"1C", x"00", x"DC", x"33", x"20", x"6D", x"6C", x"C4", x"01", x"56", x"58", x"F1", x"FE",
		x"3C", x"03", x"02", x"4D", x"50", x"63", x"4F", x"34", x"13", x"00", x"37", x"CF", x"90", x"58", x"CD", x"04",
		x"01", x"6F", x"0D", x"71", x"BF", x"0C", x"03", x"1C", x"3F", x"42", x"EF", x"A6", x"0D", x"48", x"01", x"DC",
		x"F3", x"C9", x"80", x"DC", x"38", x"00", x"EE", x"47", x"34", x"FE", x"89", x"1D", x"0A", x"F8", x"C0", x"1F",
		x"66", x"01", x"0E", x"00", x"C7", x"1F", x"FE", x"B0", x"62", x"2B", x"00", x"BB", x"BD", x"83", x"25", x"0F",
		x"74", x"00", x"BE", x"46", x"CF", x"59", x"83", x"29", x"01", x"C7", x"03", x"87", x"6D", x"87", x"25", x"00",
		x"E6", x"B0", x"F7", x"C1", x"79", x"06", x"04", x"AC", x"61", x"73", x"EC", x"8B", x"11", x"04", x"6D", x"0C",
		x"71", x"3B", x"2F", x"AC", x"00", x"DF", x"19", x"9E", x"E6", x"C0", x"2E", x"02", x"EC", x"B2", x"FF", x"0F",
		x"3E", x"00", x"0A", x"F8", x"62", x"0E", x"AC", x"1F", x"E0", x"00", x"56", x"DC", x"FF", x"A1", x"B0", x"15",
		x"00", x"7F", x"5E", x"D0", x"E8", x"81", x"E0", x"00", x"FC", x"61", x"05", x"D3", x"DE", x"D1", x"01", x"66",
		x"41", x"7F", x"23", x"9E", x"25", x"00", x"ED", x"79", x"20", x"E0", x"CE", x"76", x"00", x"E9", x"6B", x"6E",
		x"3C", x"52", x"5C", x"00", x"BF", x"1B", x"3D", x"B1", x"06", x"9C", x"03", x"3F", x"0B", x"70", x"D3", x"78",
		x"A4", x"03", x"D6", x"86", x"71", x"AC", x"65", x"0C", x"01", x"BB", x"E7", x"68", x"03", x"E2", x"C6", x"01",
		x"EB", x"37", x"86", x"D8", x"3B", x"38", x"38", x"BF", x"83", x"3D", x"F1", x"04", x"4B", x"04", x"4D", x"E1",
		x"3F", x"E3", x"C0", x"8A", x"00", x"67", x"DB", x"C1", x"5A", x"1E", x"E8", x"00", x"DD", x"CF", x"51", x"9A",
		x"C6", x"E9", x"00", x"DC", x"B3", x"E4", x"F9", x"00", x"E1", x"00", x"37", x"BF", x"C0", x"27", x"C0", x"71",
		x"00", x"AC", x"C1", x"BB", x"F9", x"0F", x"26", x"14", x"D3", x"C6", x"80", x"76", x"0F", x"53", x"00", x"CE",
		x"63", x"13", x"AC", x"B0", x"15", x"00", x"BD", x"3D", x"80", x"E0", x"5B", x"10", x"00", x"B5", x"05", x"4F",
		x"E3", x"B0", x"15", x"00", x"BF", x"A2", x"A7", x"71", x"3C", x"0B", x"02", x"37", x"BF", x"C0", x"07", x"0B",
		x"50", x"00", x"B7", x"FF", x"05", x"A2", x"C1", x"84", x"02", x"EC", x"C6", x"27", x"2C", x"63", x"19", x"07",
		x"33", x"C1", x"BE", x"21", x"B9", x"21", x"01", x"B7", x"5F", x"F0", x"32", x"80", x"5D", x"04", x"B3", x"1E",
		x"59", x"03", x"CA", x"88", x"00", x"56", x"0F", x"2F", x"28", x"6C", x"05", x"00", x"B6", x"43", x"6B", x"C8",
		x"6F", x"0B", x"10", x"37", x"6B", x"08", x"1B", x"A0", x"00", x"00", x"CF", x"02", x"B4", x"39", x"DE", x"16",
		x"00", x"D7", x"7F", x"43", x"60", x"6B", x"40", x"01", x"7E", x"1A", x"3D", x"D1", x"06", x"A4", x"00", x"4D",
		x"0F", x"4F", x"E3", x"C0", x"0A", x"00", x"3B", x"D8", x"17", x"18", x"D1", x"76", x"00", x"6F", x"87", x"A6",
		x"4D", x"80", x"05", x"01", x"5B", x"31", x"3E", x"A6", x"C0", x"12", x"00", x"67", x"03", x"3E", x"66", x"87",
		x"AD", x"08", x"76", x"1B", x"43", x"DE", x"0E", x"C6", x"10", x"F9", x"01", x"3E", x"B0", x"43", x"3B", x"00",
		x"19", x"8B", x"E7", x"13", x"E0", x"38", x"00", x"EC", x"F2", x"B3", x"00", x"95", x"15", x"00", x"59", x"43",
		x"1A", x"33", x"1E", x"29", x"00", x"9A", x"DF", x"80", x"66", x"0D", x"26", x"1C", x"56", x"58", x"1F", x"9C",
		x"67", x"09", x"00", x"37", x"16", x"B4", x"7D", x"03", x"A2", x"00", x"03", x"EE", x"BF", x"8D", x"00", x"4B",
		x"00", x"DF", x"30", x"A2", x"69", x"3C", x"52", x"00", x"56", x"AF", x"7F", x"C2", x"C1", x"06", x"04", x"56",
		x"58", x"B1", x"FF", x"83", x"05", x"01", x"76", x"83", x"F9", x"18", x"0B", x"D6", x"01", x"DF", x"92", x"A7",
		x"D1", x"80", x"A6", x"00", x"BF", x"C2", x"9E", x"D0", x"78", x"44", x"01", x"B5", x"01", x"68", x"EF", x"B0",
		x"05", x"01", x"5B", x"F1", x"0A", x"32", x"BF", x"E0", x"00", x"FC", x"82", x"09", x"56", x"AF", x"71", x"00",
		x"58", x"3F", x"86", x"BC", x"C2", x"12", x"01", x"2D", x"F1", x"3E", x"E6", x"C0", x"88", x"00", x"EC", x"60",
		x"34", x"1A", x"6F", x"C2", x"01", x"DC", x"B3", x"8C", x"B0", x"05", x"71", x"00", x"76", x"03", x"B4", x"7D",
		x"8F", x"11", x"1C", x"6B", x"F1", x"7C", x"80", x"60", x"1D", x"00", x"4D", x"F1", x"5E", x"38", x"C3", x"88",
		x"00", x"3C", x"80", x"F0", x"07", x"04", x"07", x"00", x"BD", x"07", x"04", x"80", x"05", x"00", x"00", x"C7",
		x"33", x"24", x"EF", x"01", x"E0", x"00", x"DF", x"07", x"26", x"34", x"86", x"1C", x"00", x"73", x"90", x"DB",
		x"34", x"1E", x"39", x"00", x"EB", x"87", x"21", x"8C", x"8F", x"61", x"08", x"B5", x"27", x"F8", x"60", x"6C",
		x"44", x"01", x"BF", x"F5", x"80", x"36", x"0D", x"B8", x"0E", x"FE", x"36", x"3C", x"F2", x"0D", x"08", x"07",
		x"37", x"DE", x"60", x"7A", x"62", x"C1", x"05", x"AE", x"F0", x"F0", x"65", x"70", x"01", x"81", x"00", x"AE",
		x"F0", x"F0", x"65", x"00", x"EE", x"62", x"3B", x"61", x"1A", x"A7", x"AC", x"60", x"02", x"F0", x"15", x"D2",
		x"16", x"24", x"B3", x"72", x"FB", x"32", x"27", x"1D", x"5B", x"A8", x"63", x"D2", x"16", x"00", x"EE", x"82",
		x"02", x"02", x"03", x"00", x"40", x"84", x"C4", x"A4", x"A0", x"A0", x"64", x"A0", x"02", x"43", x"00", x"40",
		x"82", x"82", x"00", x"80", x"85", x"E5", x"90", x"E0", x"84", x"A0", x"C0", x"A4", x"A4", x"40", x"40", x"A4",
		x"A0", x"40", x"80", x"44", x"A0", x"20", x"C3", x"83", x"80", x"80", x"43", x"83", x"C0", x"80", x"44", x"A0",
		x"80", x"64", x"80", x"80", x"65", x"90", x"90", x"64", x"80", x"20", x"C4", x"20", x"A0", x"60", x"E4", x"20",
		x"80", x"E0", x"15", x"75", x"90", x"70", x"10", x"F6", x"A8", x"AE", x"A8", x"50", x"50", x"AD", x"F3", x"F8",
		x"1E", x"F5", x"65", x"78", x"02", x"6A", x"F8", x"66", x"02", x"F6", x"15", x"AD", x"F7", x"F8", x"1E", x"78",
		x"01", x"F0", x"65", x"40", x"FF", x"00", x"EE", x"AD", x"6F", x"F0", x"1E", x"F3", x"65", x"86", x"00", x"80",
		x"A2", x"81", x"A2", x"82", x"A2", x"83", x"A2", x"A2", x"08", x"F3", x"55", x"A2", x"08", x"D4", x"54", x"84",
		x"64", x"84", x"05", x"24", x"B3", x"1D", x"C7", x"2A", x"1B", x"4A", x"3B", x"12", x"2C", x"02", x"02", x"02",
		x"FF", x"2D", x"1B", x"07", x"12", x"32", x"2F", x"11", x"FF", x"2A", x"1B", x"27", x"2F", x"2C", x"27", x"20",
		x"0B", x"FF", x"2A", x"1B", x"44", x"08", x"12", x"2C", x"0B", x"FF", x"30", x"1B", x"35", x"19", x"FF", x"2D",
		x"1B", x"28", x"35", x"32", x"19", x"FF", x"2C", x"1B", x"15", x"3B", x"32", x"19", x"FF", x"02", x"01", x"32",
		x"06", x"35", x"35", x"38", x"2F", x"01", x"15", x"35", x"3B", x"27", x"43", x"38", x"2F", x"2C", x"FF", x"01",
		x"0A", x"2C", x"27", x"3B", x"2B", x"2B", x"12", x"32", x"01", x"0E", x"3B", x"48", x"01", x"16", x"08", x"3F",
		x"3F", x"28", x"2F", x"FF", x"0C", x"18", x"16", x"27", x"2F", x"38", x"38", x"01", x"3B", x"01", x"19", x"2F",
		x"20", x"FF", x"0D", x"03", x"4A", x"2F", x"28", x"28", x"01", x"43", x"35", x"07", x"2F", x"11", x"FF", x"01",
		x"0A", x"08", x"07", x"28", x"35", x"32", x"19", x"2F", x"43", x"01", x"07", x"2F", x"1D", x"2C", x"01", x"38",
		x"2F", x"2C", x"FF", x"02", x"11", x"16", x"3B", x"38", x"38", x"4A", x"35", x"27", x"43", x"0D", x"FF", x"30",
		x"1B", x"07", x"35", x"FF", x"18", x"12", x"16", x"28", x"3B", x"20", x"FF", x"14", x"18", x"08", x"07", x"28",
		x"35", x"32", x"19", x"FF", x"01", x"0A", x"35", x"27", x"12", x"24", x"0D", x"01", x"07", x"35", x"15", x"03",
		x"2C", x"06", x"12", x"07", x"19", x"2B", x"08", x"07", x"FF", x"02", x"11", x"2B", x"35", x"27", x"01", x"00",
		x"32", x"06", x"12", x"16", x"00", x"01", x"15", x"20", x"01", x"06", x"3B", x"16", x"02", x"FF", x"60", x"13",
		x"24", x"B1", x"2D", x"BD", x"A8", x"04", x"F3", x"65", x"80", x"0E", x"80", x"0E", x"80", x"11", x"83", x"3E",
		x"83", x"3E", x"83", x"21", x"61", x"0A", x"62", x"05", x"82", x"03", x"81", x"33", x"A2", x"08", x"F3", x"55",
		x"63", x"2B", x"61", x"10", x"62", x"00", x"A2", x"08", x"F2", x"1E", x"F0", x"65", x"F0", x"29", x"60", x"11",
		x"24", x"B1", x"D3", x"15", x"73", x"05", x"72", x"01", x"32", x"04", x"1E", x"F6", x"00", x"EE", x"00", x"E0",
		x"68", x"AD", x"2D", x"BD", x"24", x"AF", x"2D", x"BD", x"60", x"6E", x"24", x"B1", x"00", x"EE", x"A8", x"29",
		x"60", x"10", x"D0", x"16", x"70", x"08", x"30", x"30", x"1F", x"22", x"00", x"EE", x"24", x"AF", x"68", x"9D",
		x"2D", x"BD", x"2D", x"BD", x"61", x"11", x"2F", x"1E", x"F3", x"0A", x"43", x"05", x"1F", x"48", x"43", x"08",
		x"1F", x"54", x"43", x"0A", x"1F", x"60", x"1F", x"38", x"41", x"11", x"1F", x"38", x"2F", x"1E", x"61", x"11",
		x"2F", x"1E", x"1F", x"38", x"41", x"17", x"1F", x"38", x"2F", x"1E", x"61", x"17", x"2F", x"1E", x"1F", x"38",
		x"60", x"01", x"F0", x"18", x"62", x"05", x"F2", x"15", x"2F", x"1E", x"73", x"FF", x"24", x"B3", x"33", x"00",
		x"1F", x"66", x"41", x"11", x"12", x"60", x"00", x"E0", x"64", x"02", x"65", x"0E", x"68", x"8C", x"2D", x"C3",
		x"AF", x"F5", x"F8", x"65", x"AD", x"03", x"D1", x"31", x"F0", x"0A", x"A2", x"08", x"F7", x"1E", x"77", x"01",
		x"F0", x"55", x"AD", x"03", x"D1", x"31", x"F0", x"29", x"D1", x"25", x"F6", x"18", x"47", x"04", x"1F", x"AC",
		x"71", x"05", x"AD", x"03", x"D1", x"31", x"E0", x"A1", x"1F", x"A6", x"1F", x"88", x"2D", x"55", x"A2", x"08",
		x"F3", x"65", x"81", x"43", x"82", x"53", x"52", x"00", x"1F", x"EE", x"51", x"30", x"1F", x"EE", x"81", x"00",
		x"82", x"30", x"80", x"06", x"80", x"06", x"83", x"36", x"83", x"36", x"81", x"62", x"82", x"62", x"41", x"00",
		x"1F", x"D6", x"40", x"00", x"1F", x"EE", x"42", x"00", x"1F", x"DE", x"41", x"00", x"1F", x"EE", x"43", x"00",
		x"1F", x"E6", x"42", x"00", x"1F", x"EE", x"A8", x"04", x"F3", x"55", x"24", x"A7", x"12", x"60", x"F4", x"18",
		x"2D", x"BD", x"24", x"AF", x"12", x"24", x"2B", x"0D", x"11", x"0A", x"05", x"03", x"00", x"98", x"6A", x"08",
		x"6B", x"04", x"66", x"00", x"67", x"04", x"A2", x"F7", x"FB", x"1E", x"F5", x"65", x"A2", x"F2", x"D0", x"11",
		x"22", x"D6", x"22", x"B4", x"22", x"24", x"22", x"3E", x"22", x"A2", x"22", x"52", x"22", x"6E", x"22", x"60",
		x"12", x"16", x"60", x"05", x"E0", x"A1", x"67", x"00", x"60", x"07", x"E0", x"A1", x"67", x"0C", x"60", x"08",
		x"E0", x"A1", x"67", x"08", x"60", x"09", x"E0", x"A1", x"67", x"04", x"00", x"EE", x"80", x"70", x"B2", x"42",
		x"75", x"FF", x"00", x"EE", x"74", x"01", x"00", x"EE", x"75", x"01", x"00", x"EE", x"74", x"FF", x"00", x"EE",
		x"A2", x"F7", x"7A", x"02", x"FA", x"1E", x"80", x"40", x"81", x"50", x"F1", x"55", x"00", x"EE", x"A2", x"F7",
		x"FB", x"1E", x"F1", x"65", x"A2", x"F3", x"D0", x"11", x"7B", x"02", x"00", x"EE", x"A2", x"F3", x"D4", x"51",
		x"3F", x"01", x"00", x"EE", x"54", x"80", x"12", x"EC", x"55", x"90", x"12", x"EC", x"60", x"02", x"F0", x"18",
		x"22", x"D6", x"76", x"01", x"22", x"D6", x"60", x"FF", x"61", x"FF", x"7B", x"FE", x"A2", x"F7", x"FB", x"1E",
		x"F1", x"55", x"7B", x"FE", x"A2", x"F7", x"FB", x"1E", x"F1", x"55", x"A2", x"F3", x"D4", x"51", x"12", x"B4",
		x"44", x"FF", x"12", x"EC", x"44", x"40", x"12", x"EC", x"45", x"FF", x"12", x"EC", x"45", x"20", x"12", x"EC",
		x"00", x"EE", x"C8", x"3F", x"C9", x"1F", x"60", x"07", x"80", x"97", x"3F", x"00", x"12", x"CA", x"60", x"36",
		x"80", x"87", x"3F", x"01", x"12", x"CA", x"12", x"B4", x"A2", x"F3", x"D8", x"91", x"4F", x"00", x"00", x"EE",
		x"D8", x"91", x"12", x"B4", x"A2", x"F4", x"F6", x"33", x"F2", x"65", x"60", x"37", x"63", x"00", x"F1", x"29",
		x"D0", x"35", x"70", x"05", x"F2", x"29", x"D0", x"35", x"00", x"EE", x"60", x"0F", x"F0", x"18", x"12", x"F0",
		x"E0", x"80", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0A", x"0A", x"0B", x"0A", x"0C", x"0A", x"12",
		x"05", x"43", x"38", x"50", x"60", x"00", x"85", x"00", x"C0", x"38", x"81", x"50", x"A5", x"B0", x"F1", x"1E",
		x"F0", x"55", x"60", x"00", x"85", x"00", x"C0", x"18", x"81", x"50", x"A5", x"B8", x"F1", x"1E", x"F0", x"55",
		x"60", x"00", x"A5", x"B0", x"F0", x"1E", x"F0", x"65", x"8A", x"00", x"60", x"00", x"A5", x"B8", x"F0", x"1E",
		x"F0", x"65", x"8B", x"00", x"60", x"00", x"A5", x"80", x"F0", x"1E", x"DA", x"B8", x"60", x"01", x"A5", x"C2",
		x"F0", x"55", x"60", x"07", x"A5", x"C4", x"F0", x"55", x"A5", x"C2", x"F0", x"65", x"85", x"00", x"C0", x"38",
		x"81", x"50", x"A5", x"B0", x"F1", x"1E", x"F0", x"55", x"60", x"00", x"A5", x"C1", x"F0", x"55", x"A5", x"C2",
		x"F0", x"65", x"85", x"00", x"60", x"01", x"81", x"00", x"80", x"50", x"80", x"15", x"A5", x"C6", x"F0", x"55",
		x"A5", x"C2", x"F0", x"65", x"A5", x"B0", x"F0", x"1E", x"F0", x"65", x"85", x"00", x"A5", x"C1", x"F0", x"65",
		x"A5", x"B0", x"F0", x"1E", x"F0", x"65", x"86", x"00", x"60", x"08", x"81", x"00", x"80", x"60", x"80", x"14",
		x"81", x"00", x"80", x"50", x"82", x"00", x"80", x"15", x"80", x"20", x"3F", x"00", x"12", x"DB", x"A5", x"C2",
		x"F0", x"65", x"A5", x"B0", x"F0", x"1E", x"F0", x"65", x"85", x"00", x"A5", x"C1", x"F0", x"65", x"A5", x"B0",
		x"F0", x"1E", x"F0", x"65", x"86", x"00", x"60", x"08", x"81", x"00", x"80", x"60", x"80", x"15", x"81", x"00",
		x"80", x"50", x"82", x"10", x"81", x"05", x"81", x"20", x"3F", x"00", x"12", x"D5", x"60", x"01", x"A5", x"C3",
		x"F0", x"55", x"12", x"DB", x"60", x"00", x"A5", x"C3", x"F0", x"55", x"A5", x"C1", x"F0", x"65", x"85", x"00",
		x"A5", x"C6", x"F0", x"65", x"81", x"00", x"80", x"50", x"82", x"10", x"81", x"05", x"81", x"20", x"90", x"10",
		x"6F", x"00", x"3F", x"01", x"13", x"01", x"A5", x"C1", x"F0", x"65", x"70", x"01", x"F0", x"55", x"12", x"71",
		x"A5", x"C3", x"F0", x"65", x"85", x"00", x"60", x"01", x"81", x"50", x"50", x"10", x"6F", x"01", x"3F", x"00",
		x"13", x"23", x"A5", x"C2", x"F0", x"65", x"85", x"00", x"C0", x"78", x"81", x"50", x"A5", x"B0", x"F1", x"1E",
		x"F0", x"55", x"A5", x"C3", x"F0", x"65", x"85", x"00", x"60", x"00", x"81", x"50", x"50", x"10", x"6F", x"01",
		x"90", x"10", x"6F", x"00", x"3F", x"00", x"12", x"59", x"A5", x"C2", x"F0", x"65", x"85", x"00", x"C0", x"18",
		x"81", x"50", x"A5", x"B8", x"F1", x"1E", x"F0", x"55", x"60", x"00", x"A5", x"C1", x"F0", x"55", x"A5", x"C2",
		x"F0", x"65", x"85", x"00", x"60", x"01", x"81", x"00", x"80", x"50", x"80", x"15", x"A5", x"C6", x"F0", x"55",
		x"A5", x"C2", x"F0", x"65", x"A5", x"B8", x"F0", x"1E", x"F0", x"65", x"85", x"00", x"A5", x"C1", x"F0", x"65",
		x"A5", x"B8", x"F0", x"1E", x"F0", x"65", x"86", x"00", x"60", x"08", x"81", x"00", x"80", x"60", x"80", x"14",
		x"81", x"00", x"80", x"50", x"82", x"00", x"80", x"15", x"80", x"20", x"3F", x"00", x"13", x"CB", x"A5", x"C2",
		x"F0", x"65", x"A5", x"B8", x"F0", x"1E", x"F0", x"65", x"85", x"00", x"A5", x"C1", x"F0", x"65", x"A5", x"B8",
		x"F0", x"1E", x"F0", x"65", x"86", x"00", x"60", x"08", x"81", x"00", x"80", x"60", x"80", x"15", x"81", x"00",
		x"80", x"50", x"82", x"10", x"81", x"05", x"81", x"20", x"3F", x"00", x"13", x"C5", x"60", x"01", x"A5", x"C3",
		x"F0", x"55", x"13", x"CB", x"60", x"00", x"A5", x"C3", x"F0", x"55", x"A5", x"C1", x"F0", x"65", x"85", x"00",
		x"A5", x"C6", x"F0", x"65", x"81", x"00", x"80", x"50", x"82", x"10", x"81", x"05", x"81", x"20", x"90", x"10",
		x"6F", x"00", x"3F", x"01", x"13", x"F1", x"A5", x"C1", x"F0", x"65", x"70", x"01", x"F0", x"55", x"13", x"61",
		x"A5", x"C3", x"F0", x"65", x"85", x"00", x"60", x"01", x"81", x"50", x"50", x"10", x"6F", x"01", x"3F", x"00",
		x"14", x"13", x"A5", x"C2", x"F0", x"65", x"85", x"00", x"C0", x"18", x"81", x"50", x"A5", x"B8", x"F1", x"1E",
		x"F0", x"55", x"A5", x"C3", x"F0", x"65", x"85", x"00", x"60", x"00", x"81", x"50", x"50", x"10", x"6F", x"01",
		x"90", x"10", x"6F", x"00", x"3F", x"00", x"13", x"49", x"A5", x"C2", x"F0", x"65", x"A5", x"B0", x"F0", x"1E",
		x"F0", x"65", x"8A", x"00", x"A5", x"C2", x"F0", x"65", x"A5", x"B8", x"F0", x"1E", x"F0", x"65", x"8B", x"00",
		x"60", x"00", x"A5", x"80", x"F0", x"1E", x"DA", x"B8", x"A5", x"C2", x"F0", x"65", x"85", x"00", x"A5", x"C4",
		x"F0", x"65", x"81", x"00", x"80", x"50", x"82", x"10", x"81", x"05", x"81", x"20", x"90", x"10", x"6F", x"00",
		x"3F", x"01", x"14", x"6F", x"A5", x"C2", x"F0", x"65", x"70", x"01", x"F0", x"55", x"12", x"49", x"C0", x"07",
		x"A5", x"C0", x"F0", x"55", x"A5", x"C0", x"F0", x"65", x"A5", x"B0", x"F0", x"1E", x"F0", x"65", x"8A", x"00",
		x"A5", x"C0", x"F0", x"65", x"A5", x"B8", x"F0", x"1E", x"F0", x"65", x"8B", x"00", x"A5", x"C0", x"F0", x"65",
		x"A5", x"A8", x"F0", x"1E", x"F0", x"65", x"A5", x"80", x"F0", x"1E", x"F0", x"65", x"DA", x"B8", x"60", x"0A",
		x"F0", x"15", x"A5", x"C0", x"F0", x"65", x"85", x"00", x"A5", x"C0", x"F0", x"65", x"A5", x"A8", x"F0", x"1E",
		x"F0", x"65", x"86", x"00", x"60", x"08", x"81", x"00", x"80", x"60", x"80", x"14", x"81", x"50", x"A5", x"A8",
		x"F1", x"1E", x"F0", x"55", x"A5", x"C0", x"F0", x"65", x"A5", x"A8", x"F0", x"1E", x"F0", x"65", x"85", x"00",
		x"60", x"20", x"81", x"00", x"80", x"50", x"82", x"10", x"81", x"05", x"81", x"20", x"3F", x"00", x"14", x"F1",
		x"A5", x"C0", x"F0", x"65", x"85", x"00", x"60", x"00", x"81", x"50", x"A5", x"A8", x"F1", x"1E", x"F0", x"55",
		x"A5", x"C0", x"F0", x"65", x"85", x"00", x"60", x"32", x"81", x"50", x"50", x"10", x"6F", x"01", x"90", x"10",
		x"6F", x"00", x"3F", x"00", x"14", x"6F", x"15", x"07", x"81", x"00", x"A5", x"C7", x"62", x"01", x"8E", x"25",
		x"FE", x"1E", x"F0", x"65", x"00", x"EE", x"62", x"01", x"63", x"00", x"83", x"04", x"81", x"25", x"31", x"00",
		x"15", x"1B", x"80", x"30", x"00", x"EE", x"A5", x"C7", x"FE", x"1E", x"F6", x"55", x"66", x"00", x"82", x"00",
		x"82", x"15", x"3F", x"01", x"15", x"53", x"83", x"00", x"83", x"06", x"84", x"10", x"65", x"01", x"82", x"30",
		x"82", x"45", x"3F", x"01", x"15", x"4D", x"84", x"0E", x"85", x"0E", x"15", x"3F", x"80", x"45", x"86", x"54",
		x"15", x"2F", x"F5", x"65", x"80", x"60", x"00", x"EE", x"82", x"00", x"80", x"15", x"3F", x"00", x"15", x"59",
		x"80", x"20", x"00", x"EE", x"A5", x"7D", x"F0", x"33", x"F2", x"65", x"F0", x"29", x"D3", x"45", x"73", x"06",
		x"F1", x"29", x"D3", x"45", x"73", x"06", x"F2", x"29", x"D3", x"45", x"00", x"EE", x"28", x"63", x"29", x"00",
		x"00", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"38", x"28", x"38", x"00", x"00", x"00", x"00",
		x"54", x"00", x"44", x"00", x"54", x"00", x"00", x"92", x"00", x"00", x"82", x"00", x"00", x"92", x"00", x"92",
		x"54", x"38", x"FE", x"38", x"54", x"92", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"12", x"12", x"8D", x"8D", x"20", x"A9", x"31", x"39", x"39",
		x"30", x"20", x"52", x"54", x"54", x"20", x"8E", x"8E", x"00", x"24", x"B6", x"24", x"DA", x"60", x"0F", x"E0",
		x"A1", x"12", x"24", x"60", x"0E", x"E0", x"A1", x"12", x"28", x"12", x"16", x"24", x"DA", x"12", x"2C", x"00",
		x"E0", x"12", x"2C", x"C1", x"1F", x"71", x"10", x"C2", x"0F", x"72", x"08", x"C3", x"03", x"85", x"30", x"86",
		x"10", x"87", x"20", x"88", x"30", x"48", x"00", x"77", x"01", x"48", x"01", x"77", x"FF", x"48", x"02", x"76",
		x"01", x"48", x"03", x"76", x"FF", x"A5", x"4C", x"D1", x"21", x"D6", x"71", x"64", x"F0", x"69", x"F1", x"A8",
		x"00", x"F4", x"1E", x"80", x"30", x"F0", x"55", x"74", x"01", x"A8", x"00", x"F4", x"1E", x"60", x"01", x"F0",
		x"55", x"25", x"22", x"6A", x"00", x"7A", x"00", x"F0", x"07", x"30", x"00", x"12", x"9C", x"3D", x"00", x"12",
		x"94", x"60", x"00", x"F0", x"29", x"DB", x"C5", x"3F", x"01", x"12", x"8C", x"DB", x"C5", x"25", x"22", x"F0",
		x"15", x"12", x"9C", x"FE", x"15", x"6D", x"01", x"6E", x"00", x"12", x"9C", x"80", x"E0", x"F0", x"29", x"DB",
		x"C5", x"25", x"22", x"60", x"03", x"E0", x"A1", x"63", x"00", x"60", x"06", x"E0", x"A1", x"63", x"01", x"60",
		x"07", x"E0", x"A1", x"63", x"02", x"60", x"08", x"E0", x"A1", x"63", x"03", x"43", x"00", x"72", x"FF", x"43",
		x"01", x"72", x"01", x"43", x"02", x"71", x"FF", x"43", x"03", x"71", x"01", x"A5", x"4C", x"D1", x"21", x"3F",
		x"01", x"13", x"24", x"3D", x"01", x"13", x"88", x"60", x"3F", x"81", x"02", x"60", x"1F", x"82", x"02", x"80",
		x"B0", x"80", x"17", x"3F", x"01", x"13", x"88", x"80", x"B0", x"70", x"03", x"80", x"15", x"3F", x"01", x"13",
		x"88", x"80", x"C0", x"80", x"27", x"3F", x"01", x"13", x"88", x"80", x"C0", x"70", x"04", x"80", x"25", x"3F",
		x"01", x"13", x"88", x"60", x"04", x"F0", x"18", x"CE", x"07", x"7E", x"02", x"8A", x"E4", x"A5", x"4C", x"D1",
		x"21", x"60", x"00", x"F0", x"29", x"DB", x"C5", x"80", x"E0", x"F0", x"29", x"DB", x"C5", x"60", x"30", x"F0",
		x"15", x"F0", x"07", x"30", x"00", x"13", x"1A", x"A5", x"4C", x"D1", x"21", x"93", x"50", x"13", x"3E", x"74",
		x"01", x"A8", x"00", x"F4", x"1E", x"80", x"30", x"F0", x"55", x"74", x"01", x"A8", x"00", x"F4", x"1E", x"60",
		x"00", x"F0", x"55", x"85", x"30", x"A8", x"00", x"F4", x"1E", x"F0", x"65", x"70", x"01", x"F0", x"55", x"4A",
		x"00", x"13", x"58", x"60", x"0C", x"70", x"FF", x"30", x"00", x"13", x"4E", x"7A", x"FF", x"12", x"70", x"A5",
		x"4C", x"D6", x"71", x"48", x"00", x"77", x"FF", x"48", x"01", x"77", x"01", x"48", x"02", x"76", x"FF", x"48",
		x"03", x"76", x"01", x"A8", x"00", x"F9", x"1E", x"F0", x"65", x"70", x"FF", x"F0", x"55", x"30", x"00", x"12",
		x"70", x"79", x"01", x"A8", x"00", x"F9", x"1E", x"F0", x"65", x"88", x"00", x"79", x"01", x"12", x"70", x"60",
		x"0D", x"F0", x"18", x"60", x"0B", x"E0", x"9E", x"13", x"8E", x"6B", x"01", x"6C", x"00", x"6D", x"00", x"7B",
		x"01", x"3B", x"0A", x"13", x"AA", x"6B", x"00", x"7C", x"01", x"3C", x"0A", x"13", x"AA", x"6C", x"00", x"7D",
		x"01", x"A5", x"4C", x"D6", x"71", x"48", x"00", x"77", x"FF", x"48", x"01", x"77", x"01", x"48", x"02", x"76",
		x"FF", x"48", x"03", x"76", x"01", x"A8", x"00", x"F9", x"1E", x"F0", x"65", x"70", x"FF", x"F0", x"55", x"30",
		x"00", x"13", x"98", x"99", x"40", x"13", x"DE", x"79", x"01", x"A8", x"00", x"F9", x"1E", x"F0", x"65", x"88",
		x"00", x"79", x"01", x"13", x"98", x"00", x"E0", x"66", x"11", x"67", x"09", x"68", x"2F", x"69", x"17", x"A5",
		x"52", x"D6", x"7E", x"D8", x"7E", x"77", x"FF", x"A5", x"4E", x"D6", x"71", x"D6", x"91", x"76", x"08", x"D6",
		x"71", x"D6", x"91", x"76", x"08", x"D6", x"71", x"D6", x"91", x"76", x"08", x"A5", x"50", x"D6", x"71", x"D6",
		x"91", x"A5", x"9E", x"66", x"13", x"67", x"11", x"24", x"9A", x"A5", x"AE", x"F3", x"65", x"93", x"D0", x"14",
		x"24", x"80", x"30", x"80", x"D5", x"3F", x"01", x"14", x"3A", x"14", x"44", x"92", x"C0", x"14", x"32", x"80",
		x"20", x"80", x"C5", x"3F", x"01", x"14", x"3A", x"14", x"44", x"80", x"10", x"80", x"B5", x"3F", x"00", x"14",
		x"44", x"A5", x"AE", x"83", x"D0", x"82", x"C0", x"81", x"B0", x"F3", x"55", x"A5", x"AE", x"F3", x"65", x"66",
		x"13", x"77", x"F9", x"8D", x"30", x"8C", x"20", x"8B", x"10", x"A5", x"A4", x"24", x"9A", x"C1", x"3F", x"C2",
		x"1F", x"60", x"0D", x"80", x"15", x"3F", x"00", x"14", x"7C", x"60", x"30", x"80", x"17", x"3F", x"00", x"14",
		x"7C", x"60", x"03", x"80", x"25", x"3F", x"00", x"14", x"7C", x"60", x"18", x"80", x"27", x"3F", x"00", x"14",
		x"7C", x"14", x"82", x"C3", x"0F", x"F3", x"29", x"D1", x"25", x"60", x"0F", x"E0", x"A1", x"14", x"90", x"60",
		x"0E", x"E0", x"A1", x"14", x"96", x"14", x"56", x"00", x"E0", x"24", x"B6", x"12", x"2C", x"00", x"E0", x"12",
		x"2C", x"D6", x"75", x"A5", x"AA", x"76", x"02", x"D6", x"74", x"FD", x"29", x"76", x"0A", x"D6", x"75", x"FC",
		x"29", x"76", x"05", x"D6", x"75", x"FB", x"29", x"76", x"05", x"D6", x"75", x"00", x"EE", x"A5", x"4E", x"61",
		x"00", x"62", x"00", x"66", x"1F", x"D1", x"21", x"D1", x"61", x"71", x"08", x"31", x"40", x"14", x"BE", x"A5",
		x"52", x"62", x"01", x"65", x"3F", x"D1", x"2F", x"D5", x"2F", x"72", x"0F", x"D1", x"2F", x"D5", x"2F", x"00",
		x"EE", x"61", x"0C", x"62", x"07", x"A5", x"62", x"D1", x"2A", x"A5", x"6C", x"71", x"06", x"D1", x"2A", x"A5",
		x"76", x"71", x"06", x"D1", x"2A", x"A5", x"6C", x"71", x"06", x"D1", x"2A", x"A5", x"80", x"71", x"06", x"D1",
		x"2A", x"A5", x"6C", x"71", x"06", x"D1", x"2A", x"61", x"0E", x"62", x"18", x"A5", x"8A", x"D1", x"23", x"A5",
		x"8E", x"71", x"08", x"72", x"FF", x"D1", x"24", x"71", x"09", x"72", x"FE", x"A5", x"92", x"D1", x"26", x"71",
		x"06", x"72", x"01", x"A5", x"98", x"D1", x"25", x"00", x"EE", x"6D", x"C5", x"CB", x"3F", x"8E", x"B0", x"8E",
		x"D4", x"4F", x"01", x"15", x"24", x"7B", x"01", x"6D", x"E6", x"CC", x"1F", x"8E", x"C0", x"8E", x"D4", x"4F",
		x"01", x"15", x"32", x"7C", x"01", x"6D", x"00", x"CE", x"3F", x"7E", x"40", x"FE", x"15", x"CE", x"3F", x"7E",
		x"40", x"00", x"EE", x"80", x"00", x"FF", x"00", x"FE", x"00", x"80", x"80", x"80", x"80", x"80", x"80", x"80",
		x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"1F", x"10", x"10", x"10", x"1F", x"01", x"01",
		x"01", x"01", x"1F", x"11", x"11", x"11", x"11", x"1F", x"04", x"04", x"04", x"04", x"04", x"1F", x"01", x"02",
		x"02", x"04", x"04", x"08", x"08", x"10", x"1F", x"1F", x"11", x"10", x"10", x"10", x"13", x"11", x"11", x"11",
		x"1F", x"05", x"05", x"02", x"00", x"71", x"51", x"51", x"75", x"0C", x"12", x"1E", x"14", x"12", x"09", x"14",
		x"3E", x"15", x"15", x"2A", x"00", x"77", x"44", x"24", x"14", x"77", x"00", x"57", x"52", x"72", x"52", x"57",
		x"00", x"00", x"01", x"00", x"01", x"00", x"00", x"00", x"00", x"12", x"30", x"76", x"FB", x"60", x"20", x"80",
		x"65", x"4F", x"00", x"66", x"00", x"13", x"84", x"00", x"FF", x"00", x"00", x"00", x"01", x"00", x"0C", x"0A",
		x"00", x"19", x"02", x"04", x"06", x"08", x"02", x"02", x"03", x"2C", x"00", x"0F", x"00", x"02", x"05", x"2E",
		x"08", x"00", x"00", x"02", x"05", x"00", x"00", x"00", x"00", x"6E", x"00", x"6D", x"A0", x"6A", x"08", x"69",
		x"06", x"68", x"04", x"67", x"02", x"66", x"19", x"64", x"10", x"63", x"0C", x"62", x"00", x"61", x"06", x"A2",
		x"12", x"FA", x"55", x"23", x"D4", x"60", x"40", x"F0", x"15", x"F0", x"07", x"30", x"00", x"12", x"50", x"23",
		x"D4", x"23", x"0A", x"23", x"62", x"A2", x"12", x"F5", x"65", x"22", x"AE", x"22", x"C6", x"22", x"EC", x"3F",
		x"01", x"23", x"14", x"3F", x"01", x"22", x"EC", x"3F", x"01", x"22", x"EC", x"3F", x"01", x"22", x"7C", x"4F",
		x"01", x"13", x"66", x"12", x"62", x"A2", x"12", x"F5", x"65", x"46", x"00", x"35", x"00", x"12", x"88", x"13",
		x"8C", x"E7", x"A1", x"62", x"09", x"E8", x"A1", x"62", x"04", x"E9", x"A1", x"62", x"06", x"EA", x"A1", x"62",
		x"01", x"42", x"00", x"00", x"EE", x"22", x"AE", x"81", x"20", x"23", x"9A", x"23", x"AC", x"6C", x"01", x"62",
		x"00", x"6F", x"00", x"A2", x"12", x"F5", x"55", x"A3", x"FF", x"41", x"01", x"60", x"00", x"41", x"04", x"60",
		x"13", x"41", x"06", x"60", x"0D", x"41", x"09", x"60", x"06", x"F0", x"1E", x"D3", x"47", x"00", x"EE", x"60",
		x"05", x"E0", x"9E", x"00", x"EE", x"45", x"0F", x"00", x"EE", x"65", x"0F", x"76", x"FF", x"A2", x"12", x"F5",
		x"55", x"74", x"03", x"73", x"03", x"23", x"9A", x"23", x"9A", x"23", x"9A", x"A2", x"23", x"F5", x"55", x"A4",
		x"19", x"D3", x"41", x"00", x"EE", x"A2", x"23", x"F5", x"65", x"45", x"00", x"00", x"EE", x"A4", x"19", x"D3",
		x"41", x"23", x"9A", x"6C", x"02", x"23", x"BE", x"4B", x"BB", x"13", x"0A", x"D3", x"41", x"A2", x"23", x"F5",
		x"55", x"00", x"EE", x"65", x"00", x"60", x"00", x"A2", x"17", x"F0", x"55", x"13", x"04", x"A2", x"1D", x"F5",
		x"65", x"35", x"0F", x"13", x"44", x"A4", x"1A", x"D3", x"45", x"32", x"00", x"13", x"32", x"C1", x"03", x"A2",
		x"19", x"F1", x"1E", x"F0", x"65", x"81", x"00", x"C2", x"0F", x"72", x"01", x"23", x"9A", x"A4", x"1A", x"6C",
		x"03", x"72", x"FF", x"6F", x"00", x"D3", x"45", x"A2", x"1D", x"F5", x"55", x"00", x"EE", x"C4", x"07", x"A4",
		x"1F", x"F4", x"1E", x"F0", x"65", x"83", x"00", x"A4", x"27", x"F4", x"1E", x"F0", x"65", x"84", x"00", x"A4",
		x"1A", x"D3", x"45", x"60", x"20", x"F0", x"18", x"65", x"0F", x"13", x"3E", x"65", x"00", x"13", x"3E", x"4C",
		x"01", x"12", x"02", x"4C", x"02", x"13", x"82", x"A2", x"23", x"F5", x"65", x"45", x"00", x"12", x"02", x"A4",
		x"19", x"D3", x"41", x"6F", x"00", x"D3", x"41", x"3F", x"01", x"12", x"02", x"7E", x"0A", x"60", x"40", x"F0",
		x"18", x"00", x"E0", x"12", x"4A", x"00", x"E0", x"23", x"D4", x"60", x"60", x"F0", x"18", x"13", x"94", x"6E",
		x"00", x"13", x"84", x"41", x"01", x"74", x"FF", x"41", x"04", x"73", x"FF", x"41", x"06", x"73", x"01", x"41",
		x"09", x"74", x"01", x"00", x"EE", x"44", x"00", x"74", x"01", x"43", x"00", x"73", x"01", x"43", x"38", x"73",
		x"FF", x"44", x"18", x"74", x"FF", x"00", x"EE", x"6B", x"00", x"44", x"00", x"13", x"CE", x"43", x"00", x"13",
		x"CE", x"43", x"3F", x"13", x"CE", x"44", x"1F", x"6B", x"BB", x"6F", x"00", x"00", x"EE", x"63", x"08", x"64",
		x"08", x"A2", x"29", x"FE", x"33", x"F2", x"65", x"23", x"EC", x"63", x"28", x"A2", x"29", x"F6", x"33", x"F2",
		x"65", x"23", x"F2", x"00", x"EE", x"F0", x"29", x"D3", x"45", x"73", x"06", x"F1", x"29", x"D3", x"45", x"73",
		x"06", x"F2", x"29", x"D3", x"45", x"00", x"EE", x"01", x"10", x"54", x"7C", x"6C", x"7C", x"7C", x"44", x"7C",
		x"7C", x"6C", x"7C", x"54", x"10", x"00", x"FC", x"78", x"6E", x"78", x"FC", x"00", x"3F", x"1E", x"76", x"1E",
		x"3F", x"00", x"80", x"A8", x"70", x"F8", x"70", x"A8", x"0B", x"1B", x"28", x"38", x"30", x"20", x"10", x"00",
		x"00", x"00", x"00", x"08", x"1B", x"1B", x"1B", x"18", x"04", x"A2", x"B4", x"23", x"E6", x"22", x"B6", x"70",
		x"01", x"D0", x"11", x"30", x"25", x"12", x"06", x"71", x"FF", x"D0", x"11", x"60", x"1A", x"D0", x"11", x"60",
		x"25", x"31", x"00", x"12", x"0E", x"C4", x"70", x"44", x"70", x"12", x"1C", x"C3", x"03", x"60", x"1E", x"61",
		x"03", x"22", x"5C", x"F5", x"15", x"D0", x"14", x"3F", x"01", x"12", x"3C", x"D0", x"14", x"71", x"FF", x"D0",
		x"14", x"23", x"40", x"12", x"1C", x"E7", x"A1", x"22", x"72", x"E8", x"A1", x"22", x"84", x"E9", x"A1", x"22",
		x"96", x"E2", x"9E", x"12", x"50", x"66", x"00", x"F6", x"15", x"F6", x"07", x"36", x"00", x"12", x"3C", x"D0",
		x"14", x"71", x"01", x"12", x"2A", x"A2", x"C4", x"F4", x"1E", x"66", x"00", x"43", x"01", x"66", x"04", x"43",
		x"02", x"66", x"08", x"43", x"03", x"66", x"0C", x"F6", x"1E", x"00", x"EE", x"D0", x"14", x"70", x"FF", x"23",
		x"34", x"3F", x"01", x"00", x"EE", x"D0", x"14", x"70", x"01", x"23", x"34", x"00", x"EE", x"D0", x"14", x"70",
		x"01", x"23", x"34", x"3F", x"01", x"00", x"EE", x"D0", x"14", x"70", x"FF", x"23", x"34", x"00", x"EE", x"D0",
		x"14", x"73", x"01", x"43", x"04", x"63", x"00", x"22", x"5C", x"23", x"34", x"3F", x"01", x"00", x"EE", x"D0",
		x"14", x"73", x"FF", x"43", x"FF", x"63", x"03", x"22", x"5C", x"23", x"34", x"00", x"EE", x"80", x"00", x"67",
		x"05", x"68", x"06", x"69", x"04", x"61", x"1F", x"65", x"10", x"62", x"07", x"00", x"EE", x"40", x"E0", x"00",
		x"00", x"40", x"C0", x"40", x"00", x"00", x"E0", x"40", x"00", x"40", x"60", x"40", x"00", x"40", x"40", x"60",
		x"00", x"20", x"E0", x"00", x"00", x"C0", x"40", x"40", x"00", x"00", x"E0", x"80", x"00", x"40", x"40", x"C0",
		x"00", x"00", x"E0", x"20", x"00", x"60", x"40", x"40", x"00", x"80", x"E0", x"00", x"00", x"40", x"C0", x"80",
		x"00", x"C0", x"60", x"00", x"00", x"40", x"C0", x"80", x"00", x"C0", x"60", x"00", x"00", x"80", x"C0", x"40",
		x"00", x"00", x"60", x"C0", x"00", x"80", x"C0", x"40", x"00", x"00", x"60", x"C0", x"00", x"C0", x"C0", x"00",
		x"00", x"C0", x"C0", x"00", x"00", x"C0", x"C0", x"00", x"00", x"C0", x"C0", x"00", x"00", x"40", x"40", x"40",
		x"40", x"00", x"F0", x"00", x"00", x"40", x"40", x"40", x"40", x"00", x"F0", x"00", x"00", x"D0", x"14", x"66",
		x"35", x"76", x"FF", x"36", x"00", x"13", x"38", x"00", x"EE", x"A2", x"B4", x"8C", x"10", x"3C", x"1E", x"7C",
		x"01", x"3C", x"1E", x"7C", x"01", x"3C", x"1E", x"7C", x"01", x"23", x"5E", x"4B", x"0A", x"23", x"72", x"91",
		x"C0", x"00", x"EE", x"71", x"01", x"13", x"50", x"60", x"1B", x"6B", x"00", x"D0", x"11", x"3F", x"00", x"7B",
		x"01", x"D0", x"11", x"70", x"01", x"30", x"25", x"13", x"62", x"00", x"EE", x"60", x"1B", x"D0", x"11", x"70",
		x"01", x"30", x"25", x"13", x"74", x"8E", x"10", x"8D", x"E0", x"7E", x"FF", x"60", x"1B", x"6B", x"00", x"D0",
		x"E1", x"3F", x"00", x"13", x"90", x"D0", x"E1", x"13", x"94", x"D0", x"D1", x"7B", x"01", x"70", x"01", x"30",
		x"25", x"13", x"86", x"4B", x"00", x"13", x"A6", x"7D", x"FF", x"7E", x"FF", x"3D", x"01", x"13", x"82", x"23",
		x"C0", x"3F", x"01", x"23", x"C0", x"7A", x"01", x"23", x"C0", x"80", x"A0", x"6D", x"07", x"80", x"D2", x"40",
		x"04", x"75", x"FE", x"45", x"02", x"65", x"04", x"00", x"EE", x"A7", x"00", x"F2", x"55", x"A8", x"04", x"FA",
		x"33", x"F2", x"65", x"F0", x"29", x"6D", x"32", x"6E", x"00", x"DD", x"E5", x"7D", x"05", x"F1", x"29", x"DD",
		x"E5", x"7D", x"05", x"F2", x"29", x"DD", x"E5", x"A7", x"00", x"F2", x"65", x"A2", x"B4", x"00", x"EE", x"6A",
		x"00", x"60", x"19", x"00", x"EE", x"37", x"23", x"12", x"18", x"54", x"49", x"43", x"54", x"41", x"43", x"20",
		x"62", x"79", x"20", x"44", x"61", x"76", x"69", x"64", x"20", x"57", x"49", x"4E", x"54", x"45", x"52", x"6B",
		x"00", x"6C", x"00", x"80", x"B0", x"81", x"C0", x"A3", x"E6", x"F1", x"55", x"A3", x"C4", x"FF", x"65", x"A3",
		x"B4", x"FF", x"55", x"A3", x"E6", x"F1", x"65", x"8B", x"00", x"8C", x"10", x"00", x"E0", x"6E", x"01", x"60",
		x"13", x"61", x"03", x"A3", x"9A", x"D0", x"11", x"70", x"08", x"30", x"2B", x"12", x"3E", x"60", x"13", x"71",
		x"08", x"31", x"23", x"12", x"3E", x"60", x"13", x"61", x"03", x"A3", x"9B", x"D0", x"1F", x"70", x"08", x"30",
		x"33", x"12", x"54", x"60", x"13", x"71", x"0F", x"D0", x"1A", x"70", x"08", x"30", x"33", x"12", x"60", x"23",
		x"66", x"F0", x"0A", x"81", x"00", x"A3", x"B4", x"F0", x"1E", x"F0", x"65", x"40", x"00", x"12", x"8A", x"22",
		x"7C", x"12", x"6A", x"60", x"10", x"F0", x"18", x"F0", x"15", x"F0", x"07", x"30", x"00", x"12", x"82", x"00",
		x"EE", x"60", x"02", x"8E", x"03", x"80", x"E0", x"F0", x"55", x"A3", x"D4", x"80", x"10", x"70", x"FF", x"80",
		x"04", x"F0", x"1E", x"F1", x"65", x"A3", x"AA", x"3E", x"03", x"A3", x"AF", x"D0", x"15", x"22", x"C8", x"3A",
		x"00", x"12", x"1C", x"A3", x"B4", x"61", x"00", x"62", x"00", x"63", x"01", x"F0", x"65", x"30", x"00", x"71",
		x"01", x"F3", x"1E", x"72", x"01", x"32", x"10", x"12", x"B4", x"31", x"10", x"12", x"6A", x"12", x"1C", x"6A",
		x"00", x"A3", x"B4", x"60", x"01", x"F0", x"1E", x"F8", x"65", x"69", x"00", x"89", x"04", x"23", x"44", x"89",
		x"14", x"23", x"44", x"89", x"24", x"23", x"4A", x"69", x"00", x"89", x"34", x"23", x"44", x"89", x"44", x"23",
		x"44", x"89", x"54", x"23", x"4A", x"69", x"00", x"89", x"64", x"23", x"44", x"89", x"74", x"23", x"44", x"89",
		x"84", x"23", x"4A", x"69", x"00", x"89", x"64", x"23", x"44", x"89", x"34", x"23", x"44", x"89", x"04", x"23",
		x"4A", x"69", x"00", x"89", x"74", x"23", x"44", x"89", x"44", x"23", x"44", x"89", x"14", x"23", x"4A", x"69",
		x"00", x"89", x"84", x"23", x"44", x"89", x"54", x"23", x"44", x"89", x"24", x"23", x"4A", x"69", x"00", x"89",
		x"84", x"23", x"44", x"89", x"44", x"23", x"44", x"89", x"04", x"23", x"4A", x"69", x"00", x"89", x"64", x"23",
		x"44", x"89", x"44", x"23", x"44", x"89", x"24", x"23", x"4A", x"00", x"EE", x"89", x"0E", x"89", x"0E", x"00",
		x"EE", x"49", x"15", x"13", x"54", x"49", x"3F", x"13", x"5A", x"00", x"EE", x"23", x"66", x"7B", x"01", x"13",
		x"5E", x"23", x"66", x"7C", x"01", x"23", x"66", x"6A", x"01", x"F0", x"0A", x"00", x"EE", x"63", x"05", x"64",
		x"0A", x"A3", x"AF", x"D3", x"45", x"63", x"02", x"74", x"06", x"A3", x"E6", x"FB", x"33", x"23", x"88", x"63",
		x"32", x"64", x"0A", x"A3", x"AA", x"D3", x"45", x"63", x"2F", x"74", x"06", x"A3", x"E6", x"FC", x"33", x"F2",
		x"65", x"F0", x"29", x"23", x"94", x"F1", x"29", x"23", x"94", x"F2", x"29", x"D3", x"45", x"73", x"05", x"00",
		x"EE", x"7F", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80", x"80",
		x"80", x"1C", x"22", x"22", x"22", x"1C", x"22", x"14", x"08", x"14", x"22", x"01", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"01", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"01", x"01", x"01", x"01", x"01", x"01", x"13", x"05", x"1B", x"05", x"23",
		x"05", x"13", x"0D", x"1B", x"0D", x"23", x"0D", x"13", x"15", x"1B", x"15", x"23", x"15", x"12", x"14", x"52",
		x"45", x"56", x"49", x"56", x"41", x"4C", x"53", x"54", x"55", x"44", x"49", x"4F", x"53", x"32", x"30", x"30",
		x"38", x"00", x"E0", x"6D", x"20", x"FD", x"15", x"23", x"BE", x"23", x"C6", x"6D", x"40", x"FD", x"15", x"23",
		x"BE", x"23", x"C6", x"6D", x"20", x"FD", x"15", x"23", x"BE", x"A4", x"83", x"24", x"48", x"6D", x"80", x"FD",
		x"15", x"23", x"BE", x"A4", x"83", x"24", x"48", x"A5", x"83", x"24", x"48", x"6D", x"00", x"6B", x"00", x"22",
		x"C6", x"4B", x"00", x"22", x"E4", x"4B", x"01", x"23", x"86", x"4B", x"02", x"22", x"EC", x"4B", x"03", x"23",
		x"86", x"4B", x"04", x"22", x"F4", x"4B", x"05", x"23", x"86", x"60", x"01", x"F0", x"15", x"23", x"BE", x"7D",
		x"01", x"60", x"3F", x"8C", x"D0", x"8C", x"02", x"4C", x"00", x"22", x"70", x"12", x"44", x"4B", x"00", x"22",
		x"90", x"4B", x"01", x"22", x"CC", x"4B", x"02", x"22", x"A2", x"4B", x"03", x"22", x"D4", x"4B", x"04", x"22",
		x"B4", x"4B", x"05", x"22", x"DC", x"7B", x"01", x"4B", x"06", x"6B", x"00", x"00", x"EE", x"23", x"08", x"C9",
		x"03", x"89", x"94", x"89", x"94", x"89", x"94", x"89", x"94", x"89", x"94", x"23", x"66", x"00", x"EE", x"22",
		x"FC", x"C9", x"03", x"89", x"94", x"89", x"94", x"89", x"94", x"89", x"94", x"89", x"94", x"23", x"66", x"00",
		x"EE", x"23", x"18", x"C9", x"03", x"89", x"94", x"89", x"94", x"89", x"94", x"89", x"94", x"89", x"94", x"23",
		x"66", x"00", x"EE", x"6E", x"00", x"23", x"08", x"00", x"EE", x"23", x"66", x"6E", x"00", x"22", x"FC", x"00",
		x"EE", x"23", x"66", x"6E", x"00", x"23", x"18", x"00", x"EE", x"23", x"66", x"6E", x"00", x"23", x"08", x"00",
		x"EE", x"23", x"08", x"7E", x"03", x"23", x"08", x"00", x"EE", x"22", x"FC", x"7E", x"02", x"22", x"FC", x"00",
		x"EE", x"23", x"18", x"7E", x"02", x"23", x"18", x"00", x"EE", x"6C", x"00", x"23", x"3A", x"23", x"3A", x"23",
		x"3A", x"23", x"3A", x"00", x"EE", x"6C", x"00", x"23", x"24", x"23", x"24", x"23", x"24", x"23", x"24", x"23",
		x"24", x"23", x"24", x"00", x"EE", x"6C", x"00", x"23", x"50", x"23", x"50", x"23", x"50", x"23", x"50", x"00",
		x"EE", x"A6", x"83", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"FC", x"1E", x"F1", x"65", x"A4",
		x"7C", x"D0", x"14", x"7C", x"02", x"00", x"EE", x"A9", x"83", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"FE",
		x"1E", x"FC", x"1E", x"F1", x"65", x"A4", x"7C", x"D0", x"14", x"7C", x"02", x"00", x"EE", x"AB", x"83", x"FE",
		x"1E", x"FE", x"1E", x"FE", x"1E", x"FE", x"1E", x"FC", x"1E", x"F1", x"65", x"A4", x"7C", x"D0", x"14", x"7C",
		x"02", x"00", x"EE", x"6C", x"00", x"60", x"1F", x"8A", x"D0", x"8A", x"C4", x"8A", x"02", x"8A", x"94", x"AD",
		x"83", x"FA", x"1E", x"FA", x"1E", x"F1", x"65", x"A4", x"80", x"D0", x"13", x"7C", x"01", x"3C", x"08", x"13",
		x"68", x"00", x"EE", x"60", x"1F", x"8A", x"D0", x"8A", x"02", x"8A", x"94", x"AD", x"83", x"FA", x"1E", x"FA",
		x"1E", x"F1", x"65", x"A4", x"80", x"D0", x"13", x"60", x"1F", x"8A", x"D0", x"7A", x"08", x"8A", x"02", x"8A",
		x"94", x"AD", x"83", x"FA", x"1E", x"FA", x"1E", x"F1", x"65", x"A4", x"80", x"D0", x"13", x"00", x"EE", x"A6",
		x"83", x"FD", x"1E", x"F0", x"65", x"30", x"00", x"F0", x"18", x"00", x"EE", x"F0", x"07", x"30", x"00", x"13",
		x"BE", x"00", x"EE", x"6D", x"04", x"61", x"0C", x"60", x"1C", x"62", x"12", x"A4", x"1E", x"F2", x"1E", x"D0",
		x"16", x"FD", x"15", x"23", x"BE", x"60", x"14", x"62", x"0C", x"A4", x"1E", x"F2", x"1E", x"D0", x"16", x"60",
		x"24", x"62", x"18", x"A4", x"1E", x"F2", x"1E", x"D0", x"16", x"FD", x"15", x"23", x"BE", x"60", x"0C", x"62",
		x"06", x"A4", x"1E", x"F2", x"1E", x"D0", x"16", x"60", x"2C", x"62", x"1E", x"A4", x"1E", x"F2", x"1E", x"D0",
		x"16", x"FD", x"15", x"23", x"BE", x"A4", x"1E", x"60", x"04", x"D0", x"16", x"60", x"34", x"62", x"24", x"A4",
		x"1E", x"F2", x"1E", x"D0", x"16", x"FD", x"15", x"23", x"BE", x"00", x"EE", x"00", x"00", x"0C", x"11", x"11",
		x"10", x"00", x"00", x"95", x"55", x"95", x"CD", x"00", x"00", x"53", x"55", x"55", x"33", x"40", x"40", x"44",
		x"42", x"41", x"46", x"00", x"40", x"6A", x"4A", x"4A", x"46", x"00", x"20", x"69", x"AA", x"AA", x"69", x"00",
		x"00", x"20", x"90", x"88", x"30", x"64", x"01", x"65", x"07", x"62", x"00", x"63", x"00", x"60", x"00", x"81",
		x"30", x"D0", x"11", x"71", x"08", x"F4", x"1E", x"D0", x"11", x"71", x"08", x"F4", x"1E", x"D0", x"11", x"71",
		x"08", x"F4", x"1E", x"D0", x"11", x"F4", x"1E", x"70", x"08", x"30", x"40", x"14", x"52", x"73", x"03", x"83",
		x"52", x"72", x"01", x"32", x"08", x"14", x"50", x"00", x"EE", x"60", x"B0", x"F0", x"60", x"40", x"A0", x"40",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"00", x"00", x"00", x"C6", x"00",
		x"00", x"00", x"DB", x"00", x"00", x"00", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"5F", x"06", x"00", x"00", x"FE", x"C6", x"00",
		x"00", x"D3", x"FB", x"00", x"00", x"F0", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"00", x"00", x"00", x"F6", x"00", x"00",
		x"00", x"FB", x"E0", x"00", x"00", x"F0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"00", x"00", x"00", x"C6", x"00",
		x"00", x"00", x"DB", x"00", x"00", x"00", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"06", x"00", x"00", x"00", x"C6", x"00",
		x"00", x"03", x"F1", x"00", x"00", x"30", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"00", x"00", x"00", x"C6", x"00", x"00",
		x"00", x"D9", x"00", x"00", x"00", x"E0", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2F", x"06", x"00", x"00", x"FF", x"C6", x"00",
		x"00", x"69", x"DB", x"00", x"00", x"E0", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"06", x"00", x"00", x"00", x"76", x"00", x"00",
		x"00", x"F3", x"E0", x"00", x"00", x"30", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"1F", x"07", x"0F", x"00", x"FF", x"FE", x"FC", x"7E", x"00", x"00", x"3E", x"7C",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"2F", x"1B", x"07", x"00", x"FF", x"F0", x"FB", x"1F", x"00", x"00", x"FE", x"B0",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"17", x"0F", x"00", x"00", x"FF", x"F8", x"7E", x"0F", x"00", x"0C", x"14", x"38",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"2F", x"0B", x"0F", x"00", x"FE", x"E0", x"FC", x"3F", x"00", x"00", x"7E", x"FC",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"17", x"1F", x"03", x"00", x"FF", x"F0", x"FF", x"1F", x"80", x"00", x"FE", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"0B", x"0F", x"00", x"00", x"FE", x"F8", x"7E", x"0F", x"00", x"1C", x"3E", x"00",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"17", x"17", x"0F", x"00", x"FE", x"C0", x"F8", x"3F", x"00", x"00", x"FE", x"FC",
		x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
		x"00", x"00", x"00", x"00", x"2B", x"1F", x"00", x"00", x"FF", x"E0", x"7F", x"1F", x"80", x"04", x"1C", x"3C",
		x"04", x"05", x"1B", x"05", x"1B", x"17", x"04", x"17", x"07", x"08", x"17", x"08", x"1C", x"08", x"15", x"1A",
		x"06", x"03", x"00", x"14", x"1B", x"0A", x"16", x"16", x"1A", x"0A", x"0E", x"1A", x"08", x"02", x"00", x"10",
		x"1E", x"0C", x"15", x"17", x"18", x"0B", x"08", x"19", x"0B", x"01", x"00", x"0D", x"20", x"0F", x"13", x"19",
		x"15", x"0A", x"03", x"15", x"20", x"12", x"0E", x"01", x"10", x"1A", x"01", x"0B", x"14", x"08", x"00", x"11",
		x"1F", x"14", x"0D", x"1B", x"12", x"01", x"04", x"09", x"15", x"06", x"00", x"0D", x"1D", x"16", x"0A", x"1B",
		x"15", x"03", x"06", x"08", x"18", x"05", x"01", x"09", x"1C", x"16", x"06", x"19", x"17", x"05", x"07", x"08",
		x"1B", x"05", x"04", x"05", x"1B", x"17", x"04", x"17", x"17", x"08", x"08", x"08", x"04", x"14", x"09", x"02",
		x"1A", x"18", x"1E", x"07", x"05", x"13", x"08", x"07", x"05", x"12", x"0E", x"01", x"19", x"19", x"1F", x"0A",
		x"02", x"12", x"08", x"06", x"08", x"12", x"14", x"02", x"18", x"1A", x"20", x"0C", x"00", x"10", x"09", x"05",
		x"0A", x"12", x"19", x"04", x"15", x"1B", x"00", x"0E", x"1F", x"0E", x"0B", x"03", x"0C", x"14", x"1D", x"08",
		x"00", x"0B", x"0E", x"01", x"11", x"1B", x"1D", x"11", x"0B", x"17", x"1F", x"0D", x"00", x"08", x"12", x"01",
		x"0D", x"1A", x"1B", x"12", x"08", x"18", x"1E", x"12", x"02", x"07", x"17", x"02", x"0A", x"17", x"19", x"13",
		x"1B", x"17", x"1B", x"05", x"04", x"17", x"04", x"05", x"17", x"08", x"17", x"14", x"1D", x"0A", x"06", x"04",
		x"15", x"1A", x"01", x"15", x"1B", x"09", x"0B", x"05", x"1B", x"0E", x"08", x"03", x"0E", x"1B", x"00", x"11",
		x"1E", x"0C", x"10", x"04", x"17", x"12", x"0A", x"02", x"08", x"1A", x"1F", x"0F", x"00", x"0D", x"16", x"04",
		x"10", x"14", x"0D", x"02", x"1E", x"14", x"03", x"16", x"1B", x"06", x"02", x"09", x"09", x"13", x"10", x"01",
		x"1A", x"18", x"1F", x"0A", x"01", x"12", x"07", x"06", x"04", x"0F", x"14", x"02", x"13", x"1B", x"20", x"0E",
		x"01", x"0E", x"0D", x"05", x"02", x"0A", x"18", x"03", x"0B", x"1B", x"1F", x"13", x"04", x"0A", x"12", x"05",
		x"04", x"17", x"04", x"05", x"1B", x"17", x"1B", x"05", x"08", x"14", x"08", x"08", x"15", x"19", x"1E", x"08",
		x"00", x"11", x"09", x"02", x"14", x"17", x"1B", x"0C", x"0E", x"17", x"1F", x"0B", x"00", x"0B", x"0F", x"01",
		x"10", x"1A", x"1C", x"10", x"09", x"13", x"1F", x"0E", x"02", x"06", x"15", x"02", x"0A", x"1A", x"1A", x"15",
		x"08", x"0E", x"1F", x"0F", x"08", x"02", x"05", x"18", x"1A", x"05", x"17", x"19", x"0A", x"09", x"1E", x"12",
		x"00", x"14", x"0E", x"01", x"11", x"1B", x"1C", x"09", x"0F", x"05", x"1D", x"14", x"00", x"0E", x"0C", x"1B",
		x"13", x"02", x"1D", x"0E", x"15", x"04", x"1C", x"15", x"00", x"0A", x"07", x"1A", x"16", x"05", x"1B", x"11",
		x"1B", x"05", x"04", x"05", x"04", x"17", x"1B", x"17", x"18", x"08", x"08", x"08", x"03", x"14", x"0A", x"02",
		x"19", x"19", x"1F", x"08", x"04", x"12", x"09", x"06", x"05", x"12", x"11", x"02", x"17", x"1A", x"20", x"0C",
		x"01", x"10", x"0A", x"05", x"07", x"11", x"17", x"03", x"14", x"1B", x"00", x"0D", x"20", x"0F", x"0C", x"03",
		x"0A", x"12", x"1C", x"07", x"00", x"0A", x"11", x"1B", x"0F", x"02", x"1E", x"11", x"0B", x"14", x"1F", x"0B",
		x"00", x"08", x"12", x"01", x"0D", x"1B", x"1B", x"13", x"0A", x"16", x"1F", x"0F", x"02", x"06", x"15", x"01",
		x"0A", x"19", x"19", x"14", x"07", x"17", x"1E", x"13", x"03", x"06", x"19", x"03", x"08", x"17", x"18", x"14",
		x"1B", x"05", x"04", x"05", x"1B", x"17", x"04", x"17", x"17", x"08", x"08", x"08", x"1B", x"08", x"16", x"1A",
		x"05", x"04", x"01", x"15", x"1A", x"09", x"17", x"15", x"1A", x"0A", x"11", x"1B", x"06", x"03", x"00", x"12",
		x"1D", x"0A", x"17", x"16", x"17", x"0A", x"0B", x"1A", x"07", x"02", x"00", x"10", x"1F", x"0C", x"16", x"17",
		x"15", x"0A", x"06", x"18", x"0A", x"01", x"20", x"0E", x"00", x"0E", x"14", x"19", x"13", x"08", x"02", x"14",
		x"20", x"11", x"0E", x"01", x"11", x"1B", x"02", x"0B", x"14", x"05", x"00", x"0F", x"1F", x"14", x"0D", x"1B",
		x"12", x"02", x"04", x"0A", x"17", x"04", x"01", x"0A", x"1D", x"15", x"08", x"1A", x"15", x"05", x"06", x"09",
		x"1B", x"17", x"1B", x"05", x"04", x"17", x"04", x"05", x"18", x"08", x"18", x"14", x"02", x"12", x"19", x"18",
		x"0A", x"02", x"1E", x"07", x"04", x"13", x"14", x"17", x"04", x"0E", x"17", x"19", x"11", x"01", x"20", x"0B",
		x"01", x"10", x"0F", x"18", x"08", x"0A", x"15", x"1A", x"17", x"02", x"20", x"0F", x"00", x"0D", x"09", x"18",
		x"0F", x"08", x"12", x"1A", x"01", x"08", x"1C", x"06", x"04", x"16", x"1D", x"13", x"16", x"09", x"0F", x"1B",
		x"05", x"04", x"00", x"12", x"1E", x"0A", x"18", x"16", x"1B", x"0D", x"0B", x"1A", x"0C", x"01", x"00", x"0E",
		x"1E", x"0E", x"12", x"17", x"1D", x"12", x"07", x"19", x"14", x"01", x"00", x"09", x"1B", x"12", x"0D", x"17",
		x"04", x"17", x"04", x"05", x"1B", x"17", x"1B", x"05", x"08", x"14", x"08", x"08", x"0A", x"03", x"01", x"14",
		x"1F", x"0B", x"16", x"1A", x"0B", x"05", x"04", x"10", x"11", x"05", x"00", x"11", x"20", x"11", x"10", x"1B",
		x"0F", x"02", x"03", x"0C", x"16", x"09", x"00", x"0E", x"1D", x"16", x"0A", x"1A", x"15", x"02", x"05", x"07",
		x"17", x"0E", x"00", x"0D", x"17", x"1A", x"1A", x"04", x"05", x"17", x"08", x"03", x"15", x"13", x"01", x"0A",
		x"1F", x"08", x"0E", x"01", x"11", x"1B", x"03", x"13", x"10", x"17", x"02", x"08", x"20", x"0E", x"13", x"01",
		x"0C", x"1A", x"02", x"0E", x"0A", x"18", x"03", x"07", x"1F", x"12", x"18", x"02", x"09", x"17", x"04", x"0B",
		x"04", x"05", x"1B", x"05", x"1B", x"17", x"04", x"17", x"1C", x"08", x"15", x"1A", x"06", x"03", x"00", x"14",
		x"1A", x"0A", x"0E", x"1A", x"08", x"02", x"00", x"10", x"18", x"0B", x"08", x"19", x"0B", x"01", x"00", x"0D",
		x"15", x"0A", x"03", x"15", x"0E", x"01", x"01", x"0B", x"14", x"08", x"00", x"11", x"12", x"01", x"14", x"12",
		x"15", x"06", x"00", x"0D", x"13", x"14", x"15", x"03", x"18", x"05", x"01", x"09", x"11", x"15", x"17", x"05",
		x"1B", x"05", x"04", x"05", x"10", x"15", x"17", x"08", x"09", x"02", x"1E", x"07", x"0E", x"15", x"08", x"07",
		x"0E", x"01", x"1F", x"0A", x"0C", x"15", x"08", x"06", x"14", x"02", x"0B", x"14", x"20", x"0C", x"09", x"05",
		x"19", x"04", x"0A", x"14", x"1F", x"0E", x"0B", x"03", x"1D", x"08", x"08", x"13", x"0E", x"01", x"1D", x"11",
		x"1F", x"0D", x"12", x"01", x"07", x"11", x"1B", x"12", x"1E", x"12", x"17", x"02", x"06", x"10", x"19", x"13",
		x"1B", x"17", x"1B", x"05", x"06", x"0E", x"17", x"08", x"1D", x"0A", x"15", x"1A", x"07", x"0C", x"1B", x"09",
		x"1B", x"0E", x"0E", x"1B", x"08", x"0A", x"1E", x"0C", x"17", x"12", x"08", x"1A", x"1F", x"0F", x"0B", x"08",
		x"10", x"14", x"1E", x"14", x"03", x"16", x"0F", x"07", x"09", x"13", x"1A", x"18", x"01", x"12", x"12", x"08",
		x"04", x"0F", x"13", x"1B", x"15", x"09", x"01", x"0E", x"02", x"0A", x"0B", x"1B", x"18", x"0B", x"04", x"0A",
		x"04", x"17", x"04", x"05", x"19", x"0E", x"08", x"14", x"00", x"11", x"09", x"02", x"18", x"10", x"06", x"12",
		x"00", x"0B", x"0F", x"01", x"16", x"13", x"05", x"10", x"02", x"06", x"14", x"14", x"15", x"02", x"05", x"0E",
		x"11", x"14", x"08", x"02", x"1A", x"05", x"05", x"0D", x"0E", x"13", x"0E", x"01", x"1C", x"09", x"06", x"0C",
		x"0D", x"11", x"13", x"02", x"1D", x"0E", x"06", x"0A", x"0E", x"0F", x"16", x"05", x"1B", x"11", x"07", x"09",
		x"10", x"0E", x"18", x"08", x"08", x"08", x"08", x"14", x"12", x"0E", x"04", x"12", x"09", x"06", x"13", x"16",
		x"14", x"0E", x"01", x"10", x"0A", x"05", x"0F", x"16", x"16", x"10", x"00", x"0D", x"0C", x"03", x"0A", x"15",
		x"16", x"12", x"00", x"0A", x"0F", x"02", x"07", x"13", x"00", x"08", x"15", x"13", x"12", x"01", x"05", x"10",
		x"02", x"06", x"15", x"01", x"13", x"15", x"05", x"0E", x"03", x"06", x"19", x"03", x"11", x"15", x"05", x"0B",
		x"1B", x"05", x"04", x"05", x"0F", x"15", x"17", x"08", x"1B", x"08", x"05", x"04", x"0E", x"15", x"1A", x"09",
		x"1A", x"0A", x"06", x"03", x"0C", x"14", x"1D", x"0A", x"17", x"0A", x"07", x"02", x"1F", x"0C", x"0B", x"14",
		x"15", x"0A", x"0A", x"01", x"20", x"0E", x"0A", x"13", x"13", x"08", x"20", x"11", x"0E", x"01", x"09", x"12",
		x"14", x"05", x"1F", x"14", x"08", x"11", x"12", x"02", x"17", x"04", x"1D", x"15", x"07", x"10", x"15", x"05",
		x"1B", x"17", x"1B", x"05", x"06", x"0E", x"18", x"08", x"19", x"18", x"1E", x"07", x"07", x"0C", x"14", x"17",
		x"17", x"19", x"20", x"0B", x"08", x"0A", x"0F", x"18", x"15", x"1A", x"0B", x"08", x"20", x"0F", x"09", x"18",
		x"12", x"1A", x"0E", x"07", x"04", x"16", x"1D", x"13", x"0F", x"1B", x"12", x"07", x"00", x"12", x"18", x"16",
		x"0B", x"1A", x"00", x"0E", x"16", x"09", x"12", x"17", x"07", x"19", x"00", x"09", x"18", x"0B", x"0D", x"17",
		x"04", x"17", x"04", x"05", x"19", x"0E", x"08", x"14", x"0A", x"03", x"01", x"14", x"18", x"10", x"0B", x"05",
		x"11", x"05", x"00", x"11", x"16", x"12", x"0F", x"02", x"16", x"09", x"00", x"0E", x"15", x"02", x"13", x"13",
		x"17", x"0E", x"00", x"0D", x"1A", x"04", x"08", x"03", x"15", x"13", x"01", x"0A", x"1F", x"08", x"0E", x"01",
		x"10", x"17", x"02", x"08", x"20", x"0E", x"13", x"01", x"0A", x"18", x"03", x"07", x"1F", x"12", x"18", x"02",
		x"10", x"0E", x"06", x"07", x"19", x"07", x"19", x"15", x"0D", x"0E", x"1B", x"09", x"16", x"17", x"09", x"05",
		x"0B", x"0E", x"1C", x"0C", x"12", x"18", x"0D", x"04", x"1C", x"0E", x"09", x"0C", x"0E", x"19", x"11", x"04",
		x"1B", x"0E", x"09", x"0A", x"0B", x"18", x"14", x"05", x"1A", x"0E", x"07", x"16", x"0A", x"09", x"14", x"12",
		x"1A", x"0E", x"05", x"14", x"0C", x"07", x"13", x"14", x"1A", x"0E", x"04", x"11", x"0E", x"07", x"11", x"15",
		x"1B", x"0E", x"04", x"0E", x"10", x"15", x"10", x"07", x"06", x"0C", x"1C", x"0F", x"0E", x"15", x"11", x"07",
		x"0A", x"0A", x"1D", x"10", x"0C", x"15", x"13", x"08", x"0E", x"0A", x"1C", x"12", x"0B", x"14", x"14", x"08",
		x"12", x"0B", x"0A", x"14", x"1A", x"14", x"05", x"08", x"15", x"0E", x"07", x"06", x"08", x"13", x"17", x"16",
		x"15", x"11", x"0A", x"04", x"07", x"11", x"17", x"0B", x"13", x"15", x"0D", x"04", x"06", x"10", x"18", x"0C",
		x"10", x"17", x"10", x"05", x"06", x"0E", x"19", x"0E", x"11", x"07", x"0B", x"17", x"18", x"10", x"07", x"0C",
		x"11", x"09", x"06", x"16", x"17", x"12", x"08", x"0A", x"10", x"0A", x"03", x"13", x"14", x"14", x"1A", x"0A",
		x"0E", x"0B", x"11", x"15", x"1D", x"0D", x"03", x"0F", x"0D", x"0A", x"1D", x"10", x"0D", x"15", x"12", x"08",
		x"0C", x"08", x"1A", x"14", x"09", x"13", x"15", x"09", x"0D", x"06", x"15", x"17", x"07", x"11", x"18", x"0B",
		x"10", x"17", x"10", x"05", x"19", x"0E", x"06", x"0E", x"0A", x"15", x"13", x"05", x"18", x"10", x"07", x"0C",
		x"06", x"10", x"17", x"05", x"16", x"13", x"09", x"0A", x"05", x"0C", x"1A", x"07", x"14", x"14", x"0C", x"09",
		x"08", x"07", x"11", x"14", x"1C", x"0A", x"05", x"11", x"0C", x"04", x"0E", x"13", x"1D", x"0D", x"04", x"0F",
		x"0D", x"11", x"11", x"03", x"1D", x"10", x"03", x"0D", x"0E", x"0F", x"16", x"04", x"1B", x"13", x"04", x"09",
		x"10", x"0E", x"19", x"07", x"06", x"07", x"06", x"15", x"12", x"0E", x"04", x"13", x"09", x"05", x"16", x"17",
		x"14", x"0E", x"03", x"10", x"0D", x"04", x"12", x"18", x"03", x"0E", x"16", x"10", x"11", x"03", x"0E", x"18",
		x"04", x"0E", x"16", x"12", x"14", x"04", x"0B", x"17", x"05", x"0E", x"18", x"06", x"15", x"13", x"0B", x"0A",
		x"05", x"0E", x"1A", x"08", x"13", x"15", x"0C", x"08", x"05", x"0E", x"1B", x"0B", x"11", x"15", x"0E", x"07",
		x"1B", x"0E", x"04", x"0E", x"0F", x"15", x"0F", x"07", x"19", x"10", x"03", x"0D", x"11", x"07", x"0E", x"15",
		x"15", x"12", x"02", x"0C", x"13", x"07", x"0C", x"14", x"11", x"12", x"03", x"0A", x"14", x"08", x"0B", x"14",
		x"0D", x"11", x"15", x"08", x"05", x"08", x"1A", x"14", x"0A", x"0E", x"18", x"16", x"17", x"09", x"08", x"06",
		x"0A", x"0B", x"15", x"18", x"18", x"0B", x"08", x"11", x"0C", x"07", x"12", x"18", x"19", x"0C", x"07", x"10",
		x"10", x"17", x"10", x"05", x"06", x"0E", x"19", x"0E", x"0E", x"15", x"14", x"05", x"07", x"0C", x"18", x"10",
		x"0E", x"13", x"19", x"06", x"08", x"0A", x"17", x"12", x"0F", x"12", x"1C", x"09", x"0B", x"08", x"05", x"12",
		x"11", x"11", x"0E", x"07", x"02", x"0F", x"1C", x"0D", x"12", x"12", x"02", x"0C", x"12", x"07", x"0D", x"14",
		x"13", x"14", x"05", x"08", x"16", x"09", x"0A", x"13", x"12", x"16", x"0A", x"05", x"18", x"0B", x"07", x"11",
		x"0F", x"17", x"10", x"05", x"19", x"0E", x"06", x"0E", x"15", x"07", x"0C", x"17", x"07", x"0C", x"18", x"10",
		x"19", x"0C", x"08", x"17", x"09", x"09", x"16", x"12", x"1A", x"10", x"05", x"15", x"0B", x"08", x"13", x"13",
		x"17", x"15", x"0E", x"08", x"03", x"12", x"1A", x"0B", x"13", x"18", x"11", x"09", x"02", x"0F", x"1B", x"0D",
		x"12", x"0B", x"0E", x"19", x"02", x"0C", x"1C", x"0F", x"11", x"0D", x"09", x"18", x"04", x"09", x"1B", x"13",
		x"10", x"10", x"0C", x"14", x"07", x"17", x"04", x"1A", x"03", x"1C", x"03", x"1D", x"05", x"1D", x"08", x"1B",
		x"0C", x"19", x"10", x"16", x"14", x"13", x"17", x"10", x"1A", x"0D", x"1B", x"0A", x"1B", x"08", x"19", x"06",
		x"17", x"05", x"13", x"06", x"10", x"07", x"0D", x"08", x"0A", x"0B", x"07", x"0E", x"06", x"10", x"06", x"12",
		x"08", x"15", x"0A", x"17", x"0D", x"18", x"10", x"19", x"13", x"19", x"16", x"18", x"18", x"17", x"19", x"14",
		x"10", x"19", x"0F", x"17", x"0D", x"17", x"0A", x"19", x"06", x"1A", x"06", x"16", x"09", x"13", x"09", x"11",
		x"07", x"10", x"03", x"0E", x"03", x"0B", x"08", x"0B", x"0B", x"0B", x"0C", x"0A", x"0C", x"06", x"0E", x"02",
		x"10", x"04", x"11", x"08", x"12", x"0A", x"14", x"09", x"19", x"07", x"1B", x"09", x"19", x"0D", x"17", x"0F",
		x"17", x"10", x"1A", x"12", x"1D", x"15", x"1A", x"16", x"15", x"15", x"14", x"16", x"13", x"18", x"12", x"1D",
		x"10", x"19", x"0E", x"17", x"0D", x"17", x"0B", x"17", x"08", x"17", x"05", x"19", x"02", x"19", x"03", x"17",
		x"08", x"14", x"0B", x"12", x"0E", x"11", x"10", x"10", x"11", x"10", x"14", x"0E", x"19", x"0B", x"1C", x"09",
		x"1C", x"09", x"19", x"09", x"17", x"0A", x"16", x"0A", x"14", x"09", x"13", x"07", x"11", x"04", x"0F", x"02",
		x"0B", x"03", x"09", x"06", x"09", x"09", x"09", x"0A", x"09", x"0B", x"08", x"0B", x"07", x"0B", x"07", x"0B",
		x"10", x"19", x"13", x"18", x"15", x"17", x"16", x"16", x"18", x"15", x"18", x"15", x"18", x"14", x"15", x"12",
		x"10", x"10", x"0B", x"0E", x"09", x"0C", x"08", x"0C", x"09", x"0B", x"0A", x"0A", x"0B", x"09", x"0D", x"08",
		x"10", x"06", x"14", x"04", x"1A", x"03", x"1D", x"04", x"1C", x"08", x"19", x"0B", x"15", x"0D", x"12", x"0F",
		x"10", x"10", x"0D", x"11", x"0A", x"13", x"06", x"16", x"03", x"19", x"03", x"1C", x"07", x"1C", x"0C", x"1A",
		x"A2", x"CD", x"69", x"38", x"6A", x"08", x"D9", x"A3", x"A2", x"D0", x"6B", x"00", x"6C", x"03", x"DB", x"C3",
		x"A2", x"D6", x"64", x"1D", x"65", x"1F", x"D4", x"51", x"67", x"00", x"68", x"0F", x"22", x"A2", x"22", x"AC",
		x"48", x"00", x"12", x"22", x"64", x"1E", x"65", x"1C", x"A2", x"D3", x"D4", x"53", x"6E", x"00", x"66", x"80",
		x"6D", x"04", x"ED", x"A1", x"66", x"FF", x"6D", x"05", x"ED", x"A1", x"66", x"00", x"6D", x"06", x"ED", x"A1",
		x"66", x"01", x"36", x"80", x"22", x"D8", x"A2", x"D0", x"DB", x"C3", x"CD", x"01", x"8B", x"D4", x"DB", x"C3",
		x"3F", x"00", x"12", x"92", x"A2", x"CD", x"D9", x"A3", x"CD", x"01", x"3D", x"00", x"6D", x"FF", x"79", x"FE",
		x"D9", x"A3", x"3F", x"00", x"12", x"8C", x"4E", x"00", x"12", x"2E", x"A2", x"D3", x"D4", x"53", x"45", x"00",
		x"12", x"86", x"75", x"FF", x"84", x"64", x"D4", x"53", x"3F", x"01", x"12", x"46", x"6D", x"08", x"8D", x"52",
		x"4D", x"08", x"12", x"8C", x"12", x"92", x"22", x"AC", x"78", x"FF", x"12", x"1E", x"22", x"A2", x"77", x"05",
		x"12", x"96", x"22", x"A2", x"77", x"0F", x"22", x"A2", x"6D", x"03", x"FD", x"18", x"A2", x"D3", x"D4", x"53",
		x"12", x"86", x"A2", x"F8", x"F7", x"33", x"63", x"00", x"22", x"B6", x"00", x"EE", x"A2", x"F8", x"F8", x"33",
		x"63", x"32", x"22", x"B6", x"00", x"EE", x"6D", x"1B", x"F2", x"65", x"F0", x"29", x"D3", x"D5", x"73", x"05",
		x"F1", x"29", x"D3", x"D5", x"73", x"05", x"F2", x"29", x"D3", x"D5", x"00", x"EE", x"01", x"7C", x"FE", x"7C",
		x"60", x"F0", x"60", x"40", x"E0", x"A0", x"F8", x"D4", x"6E", x"01", x"6D", x"10", x"FD", x"18", x"00", x"EE",
		x"00", x"E0", x"23", x"B6", x"60", x"07", x"E0", x"9E", x"12", x"04", x"68", x"00", x"67", x"03", x"23", x"46",
		x"22", x"4A", x"22", x"C0", x"23", x"66", x"23", x"8A", x"23", x"AC", x"F0", x"0A", x"22", x"5A", x"22", x"5A",
		x"22", x"D0", x"22", x"88", x"3A", x"00", x"12", x"1C", x"6C", x"01", x"23", x"AC", x"77", x"FF", x"23", x"AC",
		x"60", x"78", x"F0", x"15", x"F0", x"07", x"30", x"00", x"12", x"34", x"37", x"00", x"12", x"1C", x"23", x"AC",
		x"60", x"07", x"E0", x"9E", x"12", x"42", x"12", x"0A", x"00", x"FD", x"69", x"10", x"60", x"02", x"A2", x"54",
		x"D0", x"95", x"00", x"EE", x"80", x"80", x"80", x"80", x"80", x"00", x"60", x"01", x"E0", x"A1", x"12", x"68",
		x"60", x"04", x"E0", x"A1", x"12", x"72", x"00", x"EE", x"80", x"90", x"70", x"FF", x"40", x"00", x"00", x"EE",
		x"12", x"7C", x"80", x"90", x"70", x"01", x"40", x"1B", x"00", x"EE", x"12", x"7C", x"61", x"02", x"A2", x"54",
		x"D1", x"95", x"D1", x"05", x"89", x"00", x"00", x"EE", x"80", x"A0", x"70", x"FE", x"30", x"00", x"00", x"EE",
		x"80", x"B0", x"80", x"95", x"4F", x"00", x"00", x"EE", x"81", x"00", x"62", x"05", x"81", x"25", x"3F", x"00",
		x"00", x"EE", x"A2", x"BA", x"F0", x"1E", x"F0", x"65", x"8D", x"00", x"4B", x"01", x"6D", x"01", x"4B", x"1E",
		x"6D", x"FF", x"6C", x"01", x"60", x"0A", x"F0", x"18", x"00", x"EE", x"FF", x"FF", x"00", x"01", x"01", x"00",
		x"CB", x"20", x"7B", x"01", x"6A", x"04", x"6C", x"01", x"6D", x"01", x"A3", x"64", x"DA", x"B1", x"00", x"EE",
		x"80", x"A0", x"81", x"B0", x"8A", x"C4", x"8B", x"D4", x"A3", x"64", x"4B", x"01", x"6D", x"01", x"4B", x"1E",
		x"6D", x"FF", x"4A", x"3E", x"6C", x"FF", x"4A", x"00", x"6C", x"01", x"D0", x"11", x"DA", x"B1", x"4F", x"00",
		x"00", x"EE", x"80", x"A0", x"61", x"21", x"80", x"15", x"4F", x"00", x"00", x"EE", x"80", x"A0", x"81", x"B0",
		x"70", x"DE", x"71", x"FF", x"62", x"FF", x"63", x"FF", x"64", x"03", x"72", x"01", x"80", x"45", x"3F", x"00",
		x"13", x"0A", x"73", x"01", x"81", x"45", x"3F", x"00", x"13", x"12", x"80", x"20", x"81", x"30", x"80", x"24",
		x"80", x"24", x"81", x"34", x"81", x"34", x"70", x"22", x"71", x"01", x"A3", x"86", x"D0", x"13", x"7E", x"FF",
		x"60", x"00", x"8C", x"07", x"60", x"02", x"F0", x"18", x"23", x"8A", x"78", x"01", x"23", x"8A", x"3E", x"00",
		x"00", x"EE", x"23", x"66", x"00", x"EE", x"00", x"E0", x"60", x"00", x"61", x"00", x"62", x"1F", x"A3", x"64",
		x"D0", x"11", x"D0", x"21", x"70", x"01", x"30", x"3F", x"13", x"50", x"D0", x"11", x"71", x"01", x"31", x"20",
		x"13", x"5A", x"00", x"EE", x"80", x"00", x"61", x"01", x"63", x"0A", x"A3", x"86", x"60", x"22", x"62", x"07",
		x"D0", x"13", x"70", x"03", x"72", x"FF", x"32", x"00", x"13", x"70", x"71", x"03", x"73", x"FF", x"33", x"00",
		x"13", x"6C", x"6E", x"46", x"00", x"EE", x"E0", x"A0", x"E0", x"00", x"A3", x"A6", x"F8", x"33", x"F2", x"65",
		x"63", x"03", x"64", x"02", x"F0", x"29", x"D3", x"45", x"73", x"05", x"F1", x"29", x"D3", x"45", x"73", x"05",
		x"F2", x"29", x"D3", x"45", x"00", x"EE", x"00", x"00", x"00", x"00", x"00", x"00", x"60", x"14", x"61", x"02",
		x"F7", x"29", x"D0", x"15", x"00", x"EE", x"60", x"0A", x"61", x"0C", x"62", x"09", x"63", x"05", x"A3", x"CE",
		x"D0", x"15", x"F3", x"1E", x"70", x"05", x"72", x"FF", x"32", x"00", x"13", x"C0", x"00", x"EE", x"90", x"90",
		x"90", x"90", x"60", x"E0", x"90", x"E0", x"90", x"E0", x"E0", x"90", x"E0", x"90", x"90", x"20", x"20", x"20",
		x"20", x"20", x"90", x"90", x"60", x"90", x"90", x"00", x"00", x"60", x"00", x"00", x"F0", x"90", x"F0", x"80",
		x"80", x"F0", x"80", x"F0", x"10", x"F0", x"E0", x"90", x"E0", x"90", x"90", x"12", x"1A", x"4A", x"4D", x"4E",
		x"20", x"31", x"39", x"39", x"31", x"20", x"53", x"4F", x"46", x"54", x"57", x"41", x"52", x"45", x"53", x"20",
		x"80", x"80", x"FF", x"00", x"00", x"63", x"00", x"67", x"00", x"00", x"E0", x"A2", x"17", x"60", x"00", x"61",
		x"00", x"D0", x"11", x"71", x"FF", x"D0", x"11", x"71", x"01", x"70", x"08", x"30", x"40", x"12", x"26", x"71",
		x"01", x"A2", x"15", x"D0", x"12", x"70", x"FF", x"D0", x"12", x"70", x"01", x"71", x"02", x"31", x"1F", x"12",
		x"38", x"60", x"08", x"61", x"10", x"62", x"04", x"64", x"37", x"65", x"0F", x"66", x"02", x"D0", x"11", x"D4",
		x"51", x"68", x"01", x"E8", x"A1", x"62", x"02", x"68", x"02", x"E8", x"A1", x"62", x"04", x"68", x"07", x"E8",
		x"A1", x"62", x"01", x"68", x"0A", x"E8", x"A1", x"62", x"03", x"68", x"0B", x"E8", x"A1", x"66", x"02", x"68",
		x"0F", x"E8", x"A1", x"66", x"04", x"68", x"0C", x"E8", x"A1", x"66", x"01", x"68", x"0D", x"E8", x"A1", x"66",
		x"03", x"42", x"01", x"71", x"FF", x"42", x"02", x"70", x"FF", x"42", x"03", x"71", x"01", x"42", x"04", x"70",
		x"01", x"46", x"01", x"75", x"FF", x"46", x"02", x"74", x"FF", x"46", x"03", x"75", x"01", x"46", x"04", x"74",
		x"01", x"D0", x"11", x"3F", x"00", x"12", x"B4", x"D4", x"51", x"3F", x"00", x"12", x"B8", x"12", x"56", x"77",
		x"01", x"12", x"BA", x"73", x"01", x"68", x"00", x"78", x"01", x"38", x"00", x"12", x"BC", x"00", x"E0", x"60",
		x"08", x"61", x"04", x"F3", x"29", x"D0", x"15", x"60", x"34", x"F7", x"29", x"D0", x"15", x"68", x"00", x"78",
		x"01", x"38", x"00", x"12", x"D4", x"43", x"08", x"12", x"E4", x"47", x"08", x"12", x"E4", x"12", x"1E", x"12",
		x"E4", x"12", x"18", x"20", x"57", x"41", x"4C", x"4C", x"20", x"62", x"79", x"20", x"44", x"61", x"76", x"69",
		x"64", x"20", x"57", x"49", x"4E", x"54", x"45", x"52", x"20", x"A2", x"E4", x"60", x"00", x"61", x"00", x"62",
		x"1E", x"D0", x"11", x"D0", x"21", x"70", x"08", x"30", x"40", x"12", x"20", x"A2", x"DF", x"60", x"3E", x"61",
		x"01", x"D0", x"15", x"71", x"05", x"31", x"1A", x"12", x"30", x"D0", x"14", x"63", x"00", x"C4", x"0F", x"74",
		x"08", x"65", x"01", x"84", x"51", x"65", x"03", x"66", x"02", x"67", x"01", x"88", x"40", x"78", x"02", x"69",
		x"01", x"6A", x"04", x"6B", x"00", x"A2", x"DA", x"D3", x"45", x"D7", x"81", x"FC", x"0A", x"22", x"C4", x"6C",
		x"01", x"FC", x"15", x"FC", x"07", x"3C", x"00", x"12", x"62", x"A2", x"DA", x"8C", x"70", x"8D", x"80", x"E9",
		x"9E", x"12", x"7C", x"44", x"01", x"12", x"7C", x"D3", x"45", x"74", x"FE", x"D3", x"45", x"EA", x"9E", x"12",
		x"8A", x"44", x"19", x"12", x"8A", x"D3", x"45", x"74", x"02", x"D3", x"45", x"87", x"54", x"88", x"64", x"47",
		x"01", x"65", x"03", x"47", x"3D", x"65", x"FD", x"48", x"01", x"66", x"02", x"48", x"1D", x"66", x"FE", x"DC",
		x"D1", x"D7", x"81", x"37", x"01", x"12", x"5E", x"8C", x"80", x"8C", x"45", x"6D", x"00", x"9C", x"D0", x"12",
		x"BE", x"7D", x"01", x"3D", x"05", x"12", x"AC", x"FC", x"0A", x"22", x"C4", x"6B", x"00", x"12", x"5C", x"22",
		x"C4", x"7B", x"01", x"12", x"5C", x"A2", x"E5", x"FB", x"33", x"6C", x"34", x"6D", x"02", x"F2", x"65", x"F1",
		x"29", x"DC", x"D5", x"7C", x"05", x"F2", x"29", x"DC", x"D5", x"00", x"EE", x"80", x"80", x"80", x"80", x"80",
		x"E0", x"E0", x"E0", x"E0", x"E0", x"FF", x"A2", x"CC", x"6A", x"07", x"61", x"00", x"6B", x"08", x"60", x"00",
		x"D0", x"11", x"70", x"08", x"7B", x"FF", x"3B", x"00", x"12", x"0A", x"71", x"04", x"7A", x"FF", x"3A", x"00",
		x"12", x"06", x"66", x"00", x"67", x"10", x"A2", x"CD", x"60", x"20", x"61", x"1E", x"D0", x"11", x"63", x"1D",
		x"62", x"3F", x"82", x"02", x"77", x"FF", x"47", x"00", x"12", x"AA", x"FF", x"0A", x"A2", x"CB", x"D2", x"31",
		x"65", x"FF", x"C4", x"01", x"34", x"01", x"64", x"FF", x"A2", x"CD", x"6C", x"00", x"6E", x"04", x"EE", x"A1",
		x"6C", x"FF", x"6E", x"06", x"EE", x"A1", x"6C", x"01", x"D0", x"11", x"80", x"C4", x"D0", x"11", x"4F", x"01",
		x"12", x"98", x"42", x"00", x"64", x"01", x"42", x"3F", x"64", x"FF", x"43", x"00", x"65", x"01", x"43", x"1F",
		x"12", x"A4", x"A2", x"CB", x"D2", x"31", x"82", x"44", x"83", x"54", x"D2", x"31", x"3F", x"01", x"12", x"42",
		x"43", x"1E", x"12", x"98", x"6A", x"02", x"FA", x"18", x"76", x"01", x"46", x"70", x"12", x"AA", x"D2", x"31",
		x"C4", x"01", x"34", x"01", x"64", x"FF", x"C5", x"01", x"35", x"01", x"65", x"FF", x"12", x"42", x"6A", x"03",
		x"FA", x"18", x"A2", x"CB", x"D2", x"31", x"73", x"FF", x"12", x"36", x"A2", x"CB", x"D2", x"31", x"12", x"28",
		x"A2", x"CD", x"D0", x"11", x"A2", x"F0", x"F6", x"33", x"F2", x"65", x"63", x"18", x"64", x"1B", x"F0", x"29",
		x"D3", x"45", x"73", x"05", x"F1", x"29", x"D3", x"45", x"73", x"05", x"F2", x"29", x"D3", x"45", x"12", x"C8",
		x"01", x"80", x"44", x"FF"
	);
begin
   process(CLK)
   begin
      if rising_edge(CLK) then
         Q <= PROGRAM(ADDR);
      end if;
   end process;
end rtl;
